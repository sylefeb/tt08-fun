`define BASIC 1
`define SPLIT_INOUTS
/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

// for tinytapeout we target ice40, but then replace SB_IO cells
// by a custom implementation
`define ICE40 1
`define SIM_SB_IO 1

module tt_um_whynot (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // https://tinytapeout.com/specs/pinouts/

  // register reset
  reg rst_n_q;
  always @(posedge clk) begin
    rst_n_q <= rst_n;
  end

  M_main main(

    .in_ui(ui_in),
    .out_uo(uo_out),

    .inout_uio_i(uio_in),
    .inout_uio_o(uio_out),
    .inout_uio_oe(uio_oe),

    .in_run(1'b1),
    .reset(~rst_n_q),
    .clock(clk)
  );

  //              vvvvv inputs when in reset to allow PMOD external takeover
  // assign uio_oe = rst_n ? {1'b1,1'b1,main_uio_oe[3],main_uio_oe[2],1'b1,main_uio_oe[1],main_uio_oe[0],1'b1} : 8'h00;

endmodule

module M_vga_M_main_demo_vga (
out_vga_hs,
out_vga_vs,
out_active,
out_vblank,
out_vga_x,
out_vga_y,
reset,
out_clock,
clock
);
output  [0:0] out_vga_hs;
output  [0:0] out_vga_vs;
output  [0:0] out_active;
output  [0:0] out_vblank;
output  [11:0] out_vga_x;
output  [10:0] out_vga_y;
input reset;
output out_clock;
input clock;
assign out_clock = clock;

reg signed [10:0] _d_xcount;
reg signed [10:0] _q_xcount;
reg signed [9:0] _d_ycount;
reg signed [9:0] _q_ycount;
reg  [0:0] _d_active_h;
reg  [0:0] _q_active_h;
reg  [0:0] _d_active_v;
reg  [0:0] _q_active_v;
reg  [0:0] _d_vga_hs;
reg  [0:0] _q_vga_hs;
reg  [0:0] _d_vga_vs;
reg  [0:0] _q_vga_vs;
reg  [0:0] _d_active;
reg  [0:0] _q_active;
reg  [0:0] _d_vblank;
reg  [0:0] _q_vblank;
reg  [11:0] _d_vga_x;
reg  [11:0] _q_vga_x;
reg  [10:0] _d_vga_y;
reg  [10:0] _q_vga_y;
assign out_vga_hs = _q_vga_hs;
assign out_vga_vs = _q_vga_vs;
assign out_active = _q_active;
assign out_vblank = _q_vblank;
assign out_vga_x = _q_vga_x;
assign out_vga_y = _q_vga_y;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
_d_xcount = _q_xcount;
_d_ycount = _q_ycount;
_d_active_h = _q_active_h;
_d_active_v = _q_active_v;
_d_vga_hs = _q_vga_hs;
_d_vga_vs = _q_vga_vs;
_d_active = _q_active;
_d_vblank = _q_vblank;
_d_vga_x = _q_vga_x;
_d_vga_y = _q_vga_y;
// _always_pre
// __block_1
_d_active_h = _q_xcount==0 ? 1:_q_xcount==640 ? 0:_q_active_h;

_d_active_v = _q_ycount==0 ? 1:_q_ycount==480 ? 0:_q_active_v;

_d_active = _d_active_h&&_d_active_v;

_d_vga_x = _d_active_h ? _q_xcount:0;

_d_vga_y = _d_active_v ? _q_ycount:0;

_d_vga_hs = _q_xcount==-144 ? 0:_q_xcount==-49 ? 1:_q_vga_hs;

_d_vga_vs = _q_ycount==-35 ? 0:_q_ycount==-34 ? 1:_q_vga_vs;

_d_vblank = _q_ycount[9+:1];

if (_q_xcount==640) begin
// __block_2
// __block_4
_d_xcount = $signed(-159);

if (_q_ycount==480) begin
// __block_5
// __block_7
_d_ycount = $signed(-44);

// __block_8
end else begin
// __block_6
// __block_9
_d_ycount = _q_ycount+1;

// __block_10
end
// 'after'
// __block_11
// __block_12
end else begin
// __block_3
// __block_13
_d_xcount = _q_xcount+1;

// __block_14
end
// 'after'
// __block_15
// __block_16
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
_q_xcount <= (reset) ? 0 : _d_xcount;
_q_ycount <= (reset) ? 0 : _d_ycount;
_q_active_h <= (reset) ? 0 : _d_active_h;
_q_active_v <= (reset) ? 0 : _d_active_v;
_q_vga_hs <= _d_vga_hs;
_q_vga_vs <= _d_vga_vs;
_q_active <= _d_active;
_q_vblank <= _d_vblank;
_q_vga_x <= _d_vga_x;
_q_vga_y <= _d_vga_y;
end

endmodule

// ==== defines ====
`undef  _c___block_1_pid
`define _c___block_1_pid (5'(_c_doomhead[{_w_vga_vga_y[2+:5],_w_vga_vga_x[2+:5]}]))
`undef  _c___block_1_bval6
`define _c___block_1_bval6 (6'({_t___block_1_q6[0+:1],_t___block_1_p6[0+:1],_t___block_1_q6[1+:1],_t___block_1_p6[1+:1],_t___block_1_q6[2+:1],_t___block_1_p6[2+:1]}))
// ===============

module M_vga_demo_M_main_demo (
out_video_r,
out_video_g,
out_video_b,
out_video_hs,
out_video_vs,
reset,
out_clock,
clock
);
output  [1:0] out_video_r;
output  [1:0] out_video_g;
output  [1:0] out_video_b;
output  [0:0] out_video_hs;
output  [0:0] out_video_vs;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [0:0] _w_vga_vga_hs;
wire  [0:0] _w_vga_vga_vs;
wire  [0:0] _w_vga_active;
wire  [0:0] _w_vga_vblank;
wire  [11:0] _w_vga_vga_x;
wire  [10:0] _w_vga_vga_y;
reg  [23:0] _t___block_1_pal;
reg  [5:0] _t___block_1_p6;
reg  [2:0] _t___block_1_q6;
reg  [1:0] _t_video_r;
reg  [1:0] _t_video_g;
reg  [1:0] _t_video_b;
reg  [0:0] _t_video_hs;
reg  [0:0] _t_video_vs;

assign out_video_r = _t_video_r;
assign out_video_g = _t_video_g;
assign out_video_b = _t_video_b;
assign out_video_hs = _t_video_hs;
assign out_video_vs = _t_video_vs;
M_vga_M_main_demo_vga vga (
.out_vga_hs(_w_vga_vga_hs),
.out_vga_vs(_w_vga_vga_vs),
.out_active(_w_vga_active),
.out_vblank(_w_vga_vblank),
.out_vga_x(_w_vga_vga_x),
.out_vga_y(_w_vga_vga_y),
.reset(reset),
.clock(clock));



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1

_t___block_1_pal = _c_sub666[`_c___block_1_pid];

_t___block_1_p6 = {_w_vga_vga_x[0+:3],_w_vga_vga_y[0+:3]};

_t___block_1_q6 = _t___block_1_p6[0+:3]^_t___block_1_p6[3+:3];


_t_video_r = _w_vga_active ? (_t___block_1_pal[12+:6]<`_c___block_1_bval6 ? 2'b00:2'b11):0;

_t_video_g = _w_vga_active ? (_t___block_1_pal[6+:6]<`_c___block_1_bval6 ? 2'b00:2'b11):0;

_t_video_b = _w_vga_active ? (_t___block_1_pal[0+:6]<`_c___block_1_bval6 ? 2'b00:2'b11):0;

_t_video_hs = _w_vga_vga_hs;

_t_video_vs = _w_vga_vga_vs;

// __block_2
// _always_post
// pipeline stage triggers
end
// ==== wires ====
wire  [4:0] _c_doomhead[6143:0];
assign _c_doomhead[0] = 5'h00;
assign _c_doomhead[1] = 5'h00;
assign _c_doomhead[2] = 5'h00;
assign _c_doomhead[3] = 5'h00;
assign _c_doomhead[4] = 5'h00;
assign _c_doomhead[5] = 5'h00;
assign _c_doomhead[6] = 5'h00;
assign _c_doomhead[7] = 5'h00;
assign _c_doomhead[8] = 5'h05;
assign _c_doomhead[9] = 5'h02;
assign _c_doomhead[10] = 5'h02;
assign _c_doomhead[11] = 5'h02;
assign _c_doomhead[12] = 5'h04;
assign _c_doomhead[13] = 5'h06;
assign _c_doomhead[14] = 5'h06;
assign _c_doomhead[15] = 5'h06;
assign _c_doomhead[16] = 5'h06;
assign _c_doomhead[17] = 5'h06;
assign _c_doomhead[18] = 5'h04;
assign _c_doomhead[19] = 5'h02;
assign _c_doomhead[20] = 5'h02;
assign _c_doomhead[21] = 5'h05;
assign _c_doomhead[22] = 5'h00;
assign _c_doomhead[23] = 5'h00;
assign _c_doomhead[24] = 5'h00;
assign _c_doomhead[25] = 5'h00;
assign _c_doomhead[26] = 5'h00;
assign _c_doomhead[27] = 5'h00;
assign _c_doomhead[28] = 5'h00;
assign _c_doomhead[29] = 5'h00;
assign _c_doomhead[30] = 5'h00;
assign _c_doomhead[31] = 5'h00;
assign _c_doomhead[32] = 5'h00;
assign _c_doomhead[33] = 5'h00;
assign _c_doomhead[34] = 5'h00;
assign _c_doomhead[35] = 5'h00;
assign _c_doomhead[36] = 5'h00;
assign _c_doomhead[37] = 5'h00;
assign _c_doomhead[38] = 5'h03;
assign _c_doomhead[39] = 5'h02;
assign _c_doomhead[40] = 5'h0e;
assign _c_doomhead[41] = 5'h15;
assign _c_doomhead[42] = 5'h01;
assign _c_doomhead[43] = 5'h0b;
assign _c_doomhead[44] = 5'h0f;
assign _c_doomhead[45] = 5'h0c;
assign _c_doomhead[46] = 5'h0c;
assign _c_doomhead[47] = 5'h0c;
assign _c_doomhead[48] = 5'h0f;
assign _c_doomhead[49] = 5'h0b;
assign _c_doomhead[50] = 5'h07;
assign _c_doomhead[51] = 5'h06;
assign _c_doomhead[52] = 5'h02;
assign _c_doomhead[53] = 5'h0e;
assign _c_doomhead[54] = 5'h02;
assign _c_doomhead[55] = 5'h03;
assign _c_doomhead[56] = 5'h00;
assign _c_doomhead[57] = 5'h00;
assign _c_doomhead[58] = 5'h00;
assign _c_doomhead[59] = 5'h00;
assign _c_doomhead[60] = 5'h00;
assign _c_doomhead[61] = 5'h00;
assign _c_doomhead[62] = 5'h00;
assign _c_doomhead[63] = 5'h00;
assign _c_doomhead[64] = 5'h00;
assign _c_doomhead[65] = 5'h00;
assign _c_doomhead[66] = 5'h00;
assign _c_doomhead[67] = 5'h00;
assign _c_doomhead[68] = 5'h00;
assign _c_doomhead[69] = 5'h03;
assign _c_doomhead[70] = 5'h02;
assign _c_doomhead[71] = 5'h06;
assign _c_doomhead[72] = 5'h01;
assign _c_doomhead[73] = 5'h0b;
assign _c_doomhead[74] = 5'h0f;
assign _c_doomhead[75] = 5'h13;
assign _c_doomhead[76] = 5'h0c;
assign _c_doomhead[77] = 5'h0f;
assign _c_doomhead[78] = 5'h0a;
assign _c_doomhead[79] = 5'h07;
assign _c_doomhead[80] = 5'h07;
assign _c_doomhead[81] = 5'h07;
assign _c_doomhead[82] = 5'h01;
assign _c_doomhead[83] = 5'h01;
assign _c_doomhead[84] = 5'h06;
assign _c_doomhead[85] = 5'h06;
assign _c_doomhead[86] = 5'h0e;
assign _c_doomhead[87] = 5'h05;
assign _c_doomhead[88] = 5'h03;
assign _c_doomhead[89] = 5'h00;
assign _c_doomhead[90] = 5'h00;
assign _c_doomhead[91] = 5'h00;
assign _c_doomhead[92] = 5'h00;
assign _c_doomhead[93] = 5'h00;
assign _c_doomhead[94] = 5'h00;
assign _c_doomhead[95] = 5'h00;
assign _c_doomhead[96] = 5'h00;
assign _c_doomhead[97] = 5'h00;
assign _c_doomhead[98] = 5'h00;
assign _c_doomhead[99] = 5'h00;
assign _c_doomhead[100] = 5'h00;
assign _c_doomhead[101] = 5'h03;
assign _c_doomhead[102] = 5'h06;
assign _c_doomhead[103] = 5'h08;
assign _c_doomhead[104] = 5'h06;
assign _c_doomhead[105] = 5'h01;
assign _c_doomhead[106] = 5'h07;
assign _c_doomhead[107] = 5'h0a;
assign _c_doomhead[108] = 5'h08;
assign _c_doomhead[109] = 5'h0b;
assign _c_doomhead[110] = 5'h01;
assign _c_doomhead[111] = 5'h09;
assign _c_doomhead[112] = 5'h06;
assign _c_doomhead[113] = 5'h06;
assign _c_doomhead[114] = 5'h06;
assign _c_doomhead[115] = 5'h06;
assign _c_doomhead[116] = 5'h02;
assign _c_doomhead[117] = 5'h0e;
assign _c_doomhead[118] = 5'h03;
assign _c_doomhead[119] = 5'h03;
assign _c_doomhead[120] = 5'h11;
assign _c_doomhead[121] = 5'h00;
assign _c_doomhead[122] = 5'h00;
assign _c_doomhead[123] = 5'h00;
assign _c_doomhead[124] = 5'h00;
assign _c_doomhead[125] = 5'h00;
assign _c_doomhead[126] = 5'h00;
assign _c_doomhead[127] = 5'h00;
assign _c_doomhead[128] = 5'h00;
assign _c_doomhead[129] = 5'h00;
assign _c_doomhead[130] = 5'h00;
assign _c_doomhead[131] = 5'h00;
assign _c_doomhead[132] = 5'h11;
assign _c_doomhead[133] = 5'h10;
assign _c_doomhead[134] = 5'h02;
assign _c_doomhead[135] = 5'h06;
assign _c_doomhead[136] = 5'h02;
assign _c_doomhead[137] = 5'h01;
assign _c_doomhead[138] = 5'h07;
assign _c_doomhead[139] = 5'h01;
assign _c_doomhead[140] = 5'h01;
assign _c_doomhead[141] = 5'h01;
assign _c_doomhead[142] = 5'h01;
assign _c_doomhead[143] = 5'h05;
assign _c_doomhead[144] = 5'h01;
assign _c_doomhead[145] = 5'h02;
assign _c_doomhead[146] = 5'h05;
assign _c_doomhead[147] = 5'h02;
assign _c_doomhead[148] = 5'h05;
assign _c_doomhead[149] = 5'h03;
assign _c_doomhead[150] = 5'h11;
assign _c_doomhead[151] = 5'h11;
assign _c_doomhead[152] = 5'h11;
assign _c_doomhead[153] = 5'h11;
assign _c_doomhead[154] = 5'h00;
assign _c_doomhead[155] = 5'h00;
assign _c_doomhead[156] = 5'h00;
assign _c_doomhead[157] = 5'h00;
assign _c_doomhead[158] = 5'h00;
assign _c_doomhead[159] = 5'h00;
assign _c_doomhead[160] = 5'h00;
assign _c_doomhead[161] = 5'h00;
assign _c_doomhead[162] = 5'h00;
assign _c_doomhead[163] = 5'h00;
assign _c_doomhead[164] = 5'h11;
assign _c_doomhead[165] = 5'h10;
assign _c_doomhead[166] = 5'h05;
assign _c_doomhead[167] = 5'h0e;
assign _c_doomhead[168] = 5'h02;
assign _c_doomhead[169] = 5'h01;
assign _c_doomhead[170] = 5'h0e;
assign _c_doomhead[171] = 5'h07;
assign _c_doomhead[172] = 5'h04;
assign _c_doomhead[173] = 5'h04;
assign _c_doomhead[174] = 5'h01;
assign _c_doomhead[175] = 5'h04;
assign _c_doomhead[176] = 5'h05;
assign _c_doomhead[177] = 5'h04;
assign _c_doomhead[178] = 5'h05;
assign _c_doomhead[179] = 5'h10;
assign _c_doomhead[180] = 5'h02;
assign _c_doomhead[181] = 5'h11;
assign _c_doomhead[182] = 5'h03;
assign _c_doomhead[183] = 5'h03;
assign _c_doomhead[184] = 5'h10;
assign _c_doomhead[185] = 5'h11;
assign _c_doomhead[186] = 5'h00;
assign _c_doomhead[187] = 5'h00;
assign _c_doomhead[188] = 5'h00;
assign _c_doomhead[189] = 5'h00;
assign _c_doomhead[190] = 5'h00;
assign _c_doomhead[191] = 5'h00;
assign _c_doomhead[192] = 5'h00;
assign _c_doomhead[193] = 5'h00;
assign _c_doomhead[194] = 5'h00;
assign _c_doomhead[195] = 5'h00;
assign _c_doomhead[196] = 5'h11;
assign _c_doomhead[197] = 5'h05;
assign _c_doomhead[198] = 5'h05;
assign _c_doomhead[199] = 5'h06;
assign _c_doomhead[200] = 5'h06;
assign _c_doomhead[201] = 5'h0e;
assign _c_doomhead[202] = 5'h01;
assign _c_doomhead[203] = 5'h0e;
assign _c_doomhead[204] = 5'h04;
assign _c_doomhead[205] = 5'h06;
assign _c_doomhead[206] = 5'h04;
assign _c_doomhead[207] = 5'h04;
assign _c_doomhead[208] = 5'h01;
assign _c_doomhead[209] = 5'h01;
assign _c_doomhead[210] = 5'h01;
assign _c_doomhead[211] = 5'h08;
assign _c_doomhead[212] = 5'h08;
assign _c_doomhead[213] = 5'h04;
assign _c_doomhead[214] = 5'h05;
assign _c_doomhead[215] = 5'h10;
assign _c_doomhead[216] = 5'h05;
assign _c_doomhead[217] = 5'h11;
assign _c_doomhead[218] = 5'h00;
assign _c_doomhead[219] = 5'h00;
assign _c_doomhead[220] = 5'h00;
assign _c_doomhead[221] = 5'h00;
assign _c_doomhead[222] = 5'h00;
assign _c_doomhead[223] = 5'h00;
assign _c_doomhead[224] = 5'h00;
assign _c_doomhead[225] = 5'h00;
assign _c_doomhead[226] = 5'h00;
assign _c_doomhead[227] = 5'h00;
assign _c_doomhead[228] = 5'h11;
assign _c_doomhead[229] = 5'h05;
assign _c_doomhead[230] = 5'h0e;
assign _c_doomhead[231] = 5'h06;
assign _c_doomhead[232] = 5'h01;
assign _c_doomhead[233] = 5'h06;
assign _c_doomhead[234] = 5'h0e;
assign _c_doomhead[235] = 5'h09;
assign _c_doomhead[236] = 5'h0e;
assign _c_doomhead[237] = 5'h06;
assign _c_doomhead[238] = 5'h01;
assign _c_doomhead[239] = 5'h09;
assign _c_doomhead[240] = 5'h0a;
assign _c_doomhead[241] = 5'h07;
assign _c_doomhead[242] = 5'h09;
assign _c_doomhead[243] = 5'h01;
assign _c_doomhead[244] = 5'h01;
assign _c_doomhead[245] = 5'h01;
assign _c_doomhead[246] = 5'h04;
assign _c_doomhead[247] = 5'h05;
assign _c_doomhead[248] = 5'h05;
assign _c_doomhead[249] = 5'h11;
assign _c_doomhead[250] = 5'h00;
assign _c_doomhead[251] = 5'h00;
assign _c_doomhead[252] = 5'h00;
assign _c_doomhead[253] = 5'h00;
assign _c_doomhead[254] = 5'h00;
assign _c_doomhead[255] = 5'h00;
assign _c_doomhead[256] = 5'h00;
assign _c_doomhead[257] = 5'h00;
assign _c_doomhead[258] = 5'h00;
assign _c_doomhead[259] = 5'h00;
assign _c_doomhead[260] = 5'h11;
assign _c_doomhead[261] = 5'h05;
assign _c_doomhead[262] = 5'h02;
assign _c_doomhead[263] = 5'h01;
assign _c_doomhead[264] = 5'h0b;
assign _c_doomhead[265] = 5'h0a;
assign _c_doomhead[266] = 5'h09;
assign _c_doomhead[267] = 5'h09;
assign _c_doomhead[268] = 5'h0a;
assign _c_doomhead[269] = 5'h0a;
assign _c_doomhead[270] = 5'h0a;
assign _c_doomhead[271] = 5'h0a;
assign _c_doomhead[272] = 5'h0a;
assign _c_doomhead[273] = 5'h0a;
assign _c_doomhead[274] = 5'h09;
assign _c_doomhead[275] = 5'h09;
assign _c_doomhead[276] = 5'h0a;
assign _c_doomhead[277] = 5'h0b;
assign _c_doomhead[278] = 5'h01;
assign _c_doomhead[279] = 5'h0e;
assign _c_doomhead[280] = 5'h05;
assign _c_doomhead[281] = 5'h11;
assign _c_doomhead[282] = 5'h00;
assign _c_doomhead[283] = 5'h00;
assign _c_doomhead[284] = 5'h00;
assign _c_doomhead[285] = 5'h00;
assign _c_doomhead[286] = 5'h00;
assign _c_doomhead[287] = 5'h00;
assign _c_doomhead[288] = 5'h00;
assign _c_doomhead[289] = 5'h00;
assign _c_doomhead[290] = 5'h00;
assign _c_doomhead[291] = 5'h00;
assign _c_doomhead[292] = 5'h11;
assign _c_doomhead[293] = 5'h05;
assign _c_doomhead[294] = 5'h06;
assign _c_doomhead[295] = 5'h07;
assign _c_doomhead[296] = 5'h0c;
assign _c_doomhead[297] = 5'h13;
assign _c_doomhead[298] = 5'h13;
assign _c_doomhead[299] = 5'h0a;
assign _c_doomhead[300] = 5'h09;
assign _c_doomhead[301] = 5'h0b;
assign _c_doomhead[302] = 5'h0b;
assign _c_doomhead[303] = 5'h0b;
assign _c_doomhead[304] = 5'h0b;
assign _c_doomhead[305] = 5'h09;
assign _c_doomhead[306] = 5'h0a;
assign _c_doomhead[307] = 5'h13;
assign _c_doomhead[308] = 5'h13;
assign _c_doomhead[309] = 5'h0c;
assign _c_doomhead[310] = 5'h07;
assign _c_doomhead[311] = 5'h02;
assign _c_doomhead[312] = 5'h05;
assign _c_doomhead[313] = 5'h11;
assign _c_doomhead[314] = 5'h00;
assign _c_doomhead[315] = 5'h00;
assign _c_doomhead[316] = 5'h00;
assign _c_doomhead[317] = 5'h00;
assign _c_doomhead[318] = 5'h00;
assign _c_doomhead[319] = 5'h00;
assign _c_doomhead[320] = 5'h00;
assign _c_doomhead[321] = 5'h00;
assign _c_doomhead[322] = 5'h00;
assign _c_doomhead[323] = 5'h00;
assign _c_doomhead[324] = 5'h11;
assign _c_doomhead[325] = 5'h05;
assign _c_doomhead[326] = 5'h06;
assign _c_doomhead[327] = 5'h07;
assign _c_doomhead[328] = 5'h0c;
assign _c_doomhead[329] = 5'h19;
assign _c_doomhead[330] = 5'h12;
assign _c_doomhead[331] = 5'h0c;
assign _c_doomhead[332] = 5'h0f;
assign _c_doomhead[333] = 5'h09;
assign _c_doomhead[334] = 5'h01;
assign _c_doomhead[335] = 5'h01;
assign _c_doomhead[336] = 5'h09;
assign _c_doomhead[337] = 5'h0f;
assign _c_doomhead[338] = 5'h0c;
assign _c_doomhead[339] = 5'h12;
assign _c_doomhead[340] = 5'h19;
assign _c_doomhead[341] = 5'h0c;
assign _c_doomhead[342] = 5'h07;
assign _c_doomhead[343] = 5'h06;
assign _c_doomhead[344] = 5'h05;
assign _c_doomhead[345] = 5'h11;
assign _c_doomhead[346] = 5'h00;
assign _c_doomhead[347] = 5'h00;
assign _c_doomhead[348] = 5'h00;
assign _c_doomhead[349] = 5'h00;
assign _c_doomhead[350] = 5'h00;
assign _c_doomhead[351] = 5'h00;
assign _c_doomhead[352] = 5'h00;
assign _c_doomhead[353] = 5'h00;
assign _c_doomhead[354] = 5'h00;
assign _c_doomhead[355] = 5'h00;
assign _c_doomhead[356] = 5'h11;
assign _c_doomhead[357] = 5'h05;
assign _c_doomhead[358] = 5'h06;
assign _c_doomhead[359] = 5'h0a;
assign _c_doomhead[360] = 5'h12;
assign _c_doomhead[361] = 5'h16;
assign _c_doomhead[362] = 5'h16;
assign _c_doomhead[363] = 5'h12;
assign _c_doomhead[364] = 5'h12;
assign _c_doomhead[365] = 5'h0c;
assign _c_doomhead[366] = 5'h0d;
assign _c_doomhead[367] = 5'h0d;
assign _c_doomhead[368] = 5'h0c;
assign _c_doomhead[369] = 5'h12;
assign _c_doomhead[370] = 5'h12;
assign _c_doomhead[371] = 5'h16;
assign _c_doomhead[372] = 5'h16;
assign _c_doomhead[373] = 5'h12;
assign _c_doomhead[374] = 5'h0a;
assign _c_doomhead[375] = 5'h06;
assign _c_doomhead[376] = 5'h05;
assign _c_doomhead[377] = 5'h11;
assign _c_doomhead[378] = 5'h00;
assign _c_doomhead[379] = 5'h00;
assign _c_doomhead[380] = 5'h00;
assign _c_doomhead[381] = 5'h00;
assign _c_doomhead[382] = 5'h00;
assign _c_doomhead[383] = 5'h00;
assign _c_doomhead[384] = 5'h00;
assign _c_doomhead[385] = 5'h00;
assign _c_doomhead[386] = 5'h00;
assign _c_doomhead[387] = 5'h0a;
assign _c_doomhead[388] = 5'h04;
assign _c_doomhead[389] = 5'h05;
assign _c_doomhead[390] = 5'h06;
assign _c_doomhead[391] = 5'h04;
assign _c_doomhead[392] = 5'h04;
assign _c_doomhead[393] = 5'h0e;
assign _c_doomhead[394] = 5'h09;
assign _c_doomhead[395] = 5'h14;
assign _c_doomhead[396] = 5'h0a;
assign _c_doomhead[397] = 5'h06;
assign _c_doomhead[398] = 5'h0a;
assign _c_doomhead[399] = 5'h0a;
assign _c_doomhead[400] = 5'h06;
assign _c_doomhead[401] = 5'h0a;
assign _c_doomhead[402] = 5'h14;
assign _c_doomhead[403] = 5'h09;
assign _c_doomhead[404] = 5'h0e;
assign _c_doomhead[405] = 5'h04;
assign _c_doomhead[406] = 5'h04;
assign _c_doomhead[407] = 5'h06;
assign _c_doomhead[408] = 5'h05;
assign _c_doomhead[409] = 5'h04;
assign _c_doomhead[410] = 5'h0a;
assign _c_doomhead[411] = 5'h00;
assign _c_doomhead[412] = 5'h00;
assign _c_doomhead[413] = 5'h00;
assign _c_doomhead[414] = 5'h00;
assign _c_doomhead[415] = 5'h00;
assign _c_doomhead[416] = 5'h00;
assign _c_doomhead[417] = 5'h00;
assign _c_doomhead[418] = 5'h00;
assign _c_doomhead[419] = 5'h0a;
assign _c_doomhead[420] = 5'h04;
assign _c_doomhead[421] = 5'h05;
assign _c_doomhead[422] = 5'h01;
assign _c_doomhead[423] = 5'h0b;
assign _c_doomhead[424] = 5'h02;
assign _c_doomhead[425] = 5'h10;
assign _c_doomhead[426] = 5'h10;
assign _c_doomhead[427] = 5'h10;
assign _c_doomhead[428] = 5'h05;
assign _c_doomhead[429] = 5'h10;
assign _c_doomhead[430] = 5'h01;
assign _c_doomhead[431] = 5'h01;
assign _c_doomhead[432] = 5'h10;
assign _c_doomhead[433] = 5'h05;
assign _c_doomhead[434] = 5'h10;
assign _c_doomhead[435] = 5'h10;
assign _c_doomhead[436] = 5'h10;
assign _c_doomhead[437] = 5'h02;
assign _c_doomhead[438] = 5'h0b;
assign _c_doomhead[439] = 5'h01;
assign _c_doomhead[440] = 5'h05;
assign _c_doomhead[441] = 5'h04;
assign _c_doomhead[442] = 5'h0a;
assign _c_doomhead[443] = 5'h00;
assign _c_doomhead[444] = 5'h00;
assign _c_doomhead[445] = 5'h00;
assign _c_doomhead[446] = 5'h00;
assign _c_doomhead[447] = 5'h00;
assign _c_doomhead[448] = 5'h00;
assign _c_doomhead[449] = 5'h00;
assign _c_doomhead[450] = 5'h00;
assign _c_doomhead[451] = 5'h01;
assign _c_doomhead[452] = 5'h04;
assign _c_doomhead[453] = 5'h04;
assign _c_doomhead[454] = 5'h0a;
assign _c_doomhead[455] = 5'h06;
assign _c_doomhead[456] = 5'h07;
assign _c_doomhead[457] = 5'h17;
assign _c_doomhead[458] = 5'h07;
assign _c_doomhead[459] = 5'h0e;
assign _c_doomhead[460] = 5'h17;
assign _c_doomhead[461] = 5'h0e;
assign _c_doomhead[462] = 5'h0d;
assign _c_doomhead[463] = 5'h0d;
assign _c_doomhead[464] = 5'h0e;
assign _c_doomhead[465] = 5'h17;
assign _c_doomhead[466] = 5'h07;
assign _c_doomhead[467] = 5'h17;
assign _c_doomhead[468] = 5'h07;
assign _c_doomhead[469] = 5'h19;
assign _c_doomhead[470] = 5'h06;
assign _c_doomhead[471] = 5'h0a;
assign _c_doomhead[472] = 5'h04;
assign _c_doomhead[473] = 5'h04;
assign _c_doomhead[474] = 5'h01;
assign _c_doomhead[475] = 5'h00;
assign _c_doomhead[476] = 5'h00;
assign _c_doomhead[477] = 5'h00;
assign _c_doomhead[478] = 5'h00;
assign _c_doomhead[479] = 5'h00;
assign _c_doomhead[480] = 5'h00;
assign _c_doomhead[481] = 5'h00;
assign _c_doomhead[482] = 5'h00;
assign _c_doomhead[483] = 5'h04;
assign _c_doomhead[484] = 5'h02;
assign _c_doomhead[485] = 5'h08;
assign _c_doomhead[486] = 5'h0a;
assign _c_doomhead[487] = 5'h01;
assign _c_doomhead[488] = 5'h0b;
assign _c_doomhead[489] = 5'h18;
assign _c_doomhead[490] = 5'h1e;
assign _c_doomhead[491] = 5'h04;
assign _c_doomhead[492] = 5'h02;
assign _c_doomhead[493] = 5'h01;
assign _c_doomhead[494] = 5'h0c;
assign _c_doomhead[495] = 5'h12;
assign _c_doomhead[496] = 5'h01;
assign _c_doomhead[497] = 5'h02;
assign _c_doomhead[498] = 5'h04;
assign _c_doomhead[499] = 5'h1e;
assign _c_doomhead[500] = 5'h18;
assign _c_doomhead[501] = 5'h0b;
assign _c_doomhead[502] = 5'h01;
assign _c_doomhead[503] = 5'h0a;
assign _c_doomhead[504] = 5'h08;
assign _c_doomhead[505] = 5'h02;
assign _c_doomhead[506] = 5'h04;
assign _c_doomhead[507] = 5'h00;
assign _c_doomhead[508] = 5'h00;
assign _c_doomhead[509] = 5'h00;
assign _c_doomhead[510] = 5'h00;
assign _c_doomhead[511] = 5'h00;
assign _c_doomhead[512] = 5'h00;
assign _c_doomhead[513] = 5'h00;
assign _c_doomhead[514] = 5'h00;
assign _c_doomhead[515] = 5'h08;
assign _c_doomhead[516] = 5'h02;
assign _c_doomhead[517] = 5'h08;
assign _c_doomhead[518] = 5'h14;
assign _c_doomhead[519] = 5'h0d;
assign _c_doomhead[520] = 5'h0f;
assign _c_doomhead[521] = 5'h0b;
assign _c_doomhead[522] = 5'h01;
assign _c_doomhead[523] = 5'h0b;
assign _c_doomhead[524] = 5'h13;
assign _c_doomhead[525] = 5'h0d;
assign _c_doomhead[526] = 5'h12;
assign _c_doomhead[527] = 5'h18;
assign _c_doomhead[528] = 5'h0d;
assign _c_doomhead[529] = 5'h13;
assign _c_doomhead[530] = 5'h0b;
assign _c_doomhead[531] = 5'h01;
assign _c_doomhead[532] = 5'h0b;
assign _c_doomhead[533] = 5'h0f;
assign _c_doomhead[534] = 5'h0d;
assign _c_doomhead[535] = 5'h14;
assign _c_doomhead[536] = 5'h08;
assign _c_doomhead[537] = 5'h02;
assign _c_doomhead[538] = 5'h08;
assign _c_doomhead[539] = 5'h00;
assign _c_doomhead[540] = 5'h00;
assign _c_doomhead[541] = 5'h00;
assign _c_doomhead[542] = 5'h00;
assign _c_doomhead[543] = 5'h00;
assign _c_doomhead[544] = 5'h00;
assign _c_doomhead[545] = 5'h00;
assign _c_doomhead[546] = 5'h00;
assign _c_doomhead[547] = 5'h01;
assign _c_doomhead[548] = 5'h02;
assign _c_doomhead[549] = 5'h01;
assign _c_doomhead[550] = 5'h0c;
assign _c_doomhead[551] = 5'h14;
assign _c_doomhead[552] = 5'h19;
assign _c_doomhead[553] = 5'h14;
assign _c_doomhead[554] = 5'h13;
assign _c_doomhead[555] = 5'h12;
assign _c_doomhead[556] = 5'h16;
assign _c_doomhead[557] = 5'h12;
assign _c_doomhead[558] = 5'h12;
assign _c_doomhead[559] = 5'h18;
assign _c_doomhead[560] = 5'h12;
assign _c_doomhead[561] = 5'h16;
assign _c_doomhead[562] = 5'h12;
assign _c_doomhead[563] = 5'h13;
assign _c_doomhead[564] = 5'h14;
assign _c_doomhead[565] = 5'h19;
assign _c_doomhead[566] = 5'h14;
assign _c_doomhead[567] = 5'h0c;
assign _c_doomhead[568] = 5'h01;
assign _c_doomhead[569] = 5'h02;
assign _c_doomhead[570] = 5'h01;
assign _c_doomhead[571] = 5'h00;
assign _c_doomhead[572] = 5'h00;
assign _c_doomhead[573] = 5'h00;
assign _c_doomhead[574] = 5'h00;
assign _c_doomhead[575] = 5'h00;
assign _c_doomhead[576] = 5'h00;
assign _c_doomhead[577] = 5'h00;
assign _c_doomhead[578] = 5'h00;
assign _c_doomhead[579] = 5'h00;
assign _c_doomhead[580] = 5'h02;
assign _c_doomhead[581] = 5'h08;
assign _c_doomhead[582] = 5'h09;
assign _c_doomhead[583] = 5'h0b;
assign _c_doomhead[584] = 5'h0f;
assign _c_doomhead[585] = 5'h0d;
assign _c_doomhead[586] = 5'h12;
assign _c_doomhead[587] = 5'h16;
assign _c_doomhead[588] = 5'h14;
assign _c_doomhead[589] = 5'h0d;
assign _c_doomhead[590] = 5'h18;
assign _c_doomhead[591] = 5'h16;
assign _c_doomhead[592] = 5'h0d;
assign _c_doomhead[593] = 5'h14;
assign _c_doomhead[594] = 5'h16;
assign _c_doomhead[595] = 5'h12;
assign _c_doomhead[596] = 5'h0d;
assign _c_doomhead[597] = 5'h0f;
assign _c_doomhead[598] = 5'h0b;
assign _c_doomhead[599] = 5'h09;
assign _c_doomhead[600] = 5'h08;
assign _c_doomhead[601] = 5'h02;
assign _c_doomhead[602] = 5'h00;
assign _c_doomhead[603] = 5'h00;
assign _c_doomhead[604] = 5'h00;
assign _c_doomhead[605] = 5'h00;
assign _c_doomhead[606] = 5'h00;
assign _c_doomhead[607] = 5'h00;
assign _c_doomhead[608] = 5'h00;
assign _c_doomhead[609] = 5'h00;
assign _c_doomhead[610] = 5'h00;
assign _c_doomhead[611] = 5'h00;
assign _c_doomhead[612] = 5'h02;
assign _c_doomhead[613] = 5'h06;
assign _c_doomhead[614] = 5'h07;
assign _c_doomhead[615] = 5'h09;
assign _c_doomhead[616] = 5'h0f;
assign _c_doomhead[617] = 5'h19;
assign _c_doomhead[618] = 5'h18;
assign _c_doomhead[619] = 5'h0d;
assign _c_doomhead[620] = 5'h0b;
assign _c_doomhead[621] = 5'h07;
assign _c_doomhead[622] = 5'h00;
assign _c_doomhead[623] = 5'h00;
assign _c_doomhead[624] = 5'h07;
assign _c_doomhead[625] = 5'h0b;
assign _c_doomhead[626] = 5'h0d;
assign _c_doomhead[627] = 5'h18;
assign _c_doomhead[628] = 5'h19;
assign _c_doomhead[629] = 5'h0f;
assign _c_doomhead[630] = 5'h09;
assign _c_doomhead[631] = 5'h07;
assign _c_doomhead[632] = 5'h06;
assign _c_doomhead[633] = 5'h02;
assign _c_doomhead[634] = 5'h00;
assign _c_doomhead[635] = 5'h00;
assign _c_doomhead[636] = 5'h00;
assign _c_doomhead[637] = 5'h00;
assign _c_doomhead[638] = 5'h00;
assign _c_doomhead[639] = 5'h00;
assign _c_doomhead[640] = 5'h00;
assign _c_doomhead[641] = 5'h00;
assign _c_doomhead[642] = 5'h00;
assign _c_doomhead[643] = 5'h00;
assign _c_doomhead[644] = 5'h00;
assign _c_doomhead[645] = 5'h06;
assign _c_doomhead[646] = 5'h0a;
assign _c_doomhead[647] = 5'h07;
assign _c_doomhead[648] = 5'h0d;
assign _c_doomhead[649] = 5'h16;
assign _c_doomhead[650] = 5'h12;
assign _c_doomhead[651] = 5'h0f;
assign _c_doomhead[652] = 5'h0e;
assign _c_doomhead[653] = 5'h06;
assign _c_doomhead[654] = 5'h08;
assign _c_doomhead[655] = 5'h08;
assign _c_doomhead[656] = 5'h06;
assign _c_doomhead[657] = 5'h0e;
assign _c_doomhead[658] = 5'h0f;
assign _c_doomhead[659] = 5'h12;
assign _c_doomhead[660] = 5'h16;
assign _c_doomhead[661] = 5'h0d;
assign _c_doomhead[662] = 5'h07;
assign _c_doomhead[663] = 5'h0a;
assign _c_doomhead[664] = 5'h06;
assign _c_doomhead[665] = 5'h00;
assign _c_doomhead[666] = 5'h00;
assign _c_doomhead[667] = 5'h00;
assign _c_doomhead[668] = 5'h00;
assign _c_doomhead[669] = 5'h00;
assign _c_doomhead[670] = 5'h00;
assign _c_doomhead[671] = 5'h00;
assign _c_doomhead[672] = 5'h00;
assign _c_doomhead[673] = 5'h00;
assign _c_doomhead[674] = 5'h00;
assign _c_doomhead[675] = 5'h00;
assign _c_doomhead[676] = 5'h00;
assign _c_doomhead[677] = 5'h02;
assign _c_doomhead[678] = 5'h13;
assign _c_doomhead[679] = 5'h07;
assign _c_doomhead[680] = 5'h12;
assign _c_doomhead[681] = 5'h18;
assign _c_doomhead[682] = 5'h0c;
assign _c_doomhead[683] = 5'h0c;
assign _c_doomhead[684] = 5'h0d;
assign _c_doomhead[685] = 5'h0f;
assign _c_doomhead[686] = 5'h09;
assign _c_doomhead[687] = 5'h09;
assign _c_doomhead[688] = 5'h0f;
assign _c_doomhead[689] = 5'h0d;
assign _c_doomhead[690] = 5'h0c;
assign _c_doomhead[691] = 5'h0c;
assign _c_doomhead[692] = 5'h18;
assign _c_doomhead[693] = 5'h12;
assign _c_doomhead[694] = 5'h07;
assign _c_doomhead[695] = 5'h13;
assign _c_doomhead[696] = 5'h02;
assign _c_doomhead[697] = 5'h00;
assign _c_doomhead[698] = 5'h00;
assign _c_doomhead[699] = 5'h00;
assign _c_doomhead[700] = 5'h00;
assign _c_doomhead[701] = 5'h00;
assign _c_doomhead[702] = 5'h00;
assign _c_doomhead[703] = 5'h00;
assign _c_doomhead[704] = 5'h00;
assign _c_doomhead[705] = 5'h00;
assign _c_doomhead[706] = 5'h00;
assign _c_doomhead[707] = 5'h00;
assign _c_doomhead[708] = 5'h00;
assign _c_doomhead[709] = 5'h0e;
assign _c_doomhead[710] = 5'h0b;
assign _c_doomhead[711] = 5'h09;
assign _c_doomhead[712] = 5'h0d;
assign _c_doomhead[713] = 5'h12;
assign _c_doomhead[714] = 5'h0c;
assign _c_doomhead[715] = 5'h0d;
assign _c_doomhead[716] = 5'h18;
assign _c_doomhead[717] = 5'h16;
assign _c_doomhead[718] = 5'h14;
assign _c_doomhead[719] = 5'h14;
assign _c_doomhead[720] = 5'h16;
assign _c_doomhead[721] = 5'h18;
assign _c_doomhead[722] = 5'h0d;
assign _c_doomhead[723] = 5'h0c;
assign _c_doomhead[724] = 5'h12;
assign _c_doomhead[725] = 5'h0d;
assign _c_doomhead[726] = 5'h09;
assign _c_doomhead[727] = 5'h0b;
assign _c_doomhead[728] = 5'h0e;
assign _c_doomhead[729] = 5'h00;
assign _c_doomhead[730] = 5'h00;
assign _c_doomhead[731] = 5'h00;
assign _c_doomhead[732] = 5'h00;
assign _c_doomhead[733] = 5'h00;
assign _c_doomhead[734] = 5'h00;
assign _c_doomhead[735] = 5'h00;
assign _c_doomhead[736] = 5'h00;
assign _c_doomhead[737] = 5'h00;
assign _c_doomhead[738] = 5'h00;
assign _c_doomhead[739] = 5'h00;
assign _c_doomhead[740] = 5'h00;
assign _c_doomhead[741] = 5'h00;
assign _c_doomhead[742] = 5'h08;
assign _c_doomhead[743] = 5'h0b;
assign _c_doomhead[744] = 5'h13;
assign _c_doomhead[745] = 5'h0d;
assign _c_doomhead[746] = 5'h01;
assign _c_doomhead[747] = 5'h06;
assign _c_doomhead[748] = 5'h1f;
assign _c_doomhead[749] = 5'h1f;
assign _c_doomhead[750] = 5'h1f;
assign _c_doomhead[751] = 5'h1f;
assign _c_doomhead[752] = 5'h1f;
assign _c_doomhead[753] = 5'h1f;
assign _c_doomhead[754] = 5'h06;
assign _c_doomhead[755] = 5'h01;
assign _c_doomhead[756] = 5'h0d;
assign _c_doomhead[757] = 5'h13;
assign _c_doomhead[758] = 5'h0b;
assign _c_doomhead[759] = 5'h08;
assign _c_doomhead[760] = 5'h00;
assign _c_doomhead[761] = 5'h00;
assign _c_doomhead[762] = 5'h00;
assign _c_doomhead[763] = 5'h00;
assign _c_doomhead[764] = 5'h00;
assign _c_doomhead[765] = 5'h00;
assign _c_doomhead[766] = 5'h00;
assign _c_doomhead[767] = 5'h00;
assign _c_doomhead[768] = 5'h00;
assign _c_doomhead[769] = 5'h00;
assign _c_doomhead[770] = 5'h00;
assign _c_doomhead[771] = 5'h00;
assign _c_doomhead[772] = 5'h00;
assign _c_doomhead[773] = 5'h00;
assign _c_doomhead[774] = 5'h0e;
assign _c_doomhead[775] = 5'h01;
assign _c_doomhead[776] = 5'h0a;
assign _c_doomhead[777] = 5'h13;
assign _c_doomhead[778] = 5'h13;
assign _c_doomhead[779] = 5'h13;
assign _c_doomhead[780] = 5'h0d;
assign _c_doomhead[781] = 5'h12;
assign _c_doomhead[782] = 5'h12;
assign _c_doomhead[783] = 5'h12;
assign _c_doomhead[784] = 5'h12;
assign _c_doomhead[785] = 5'h0d;
assign _c_doomhead[786] = 5'h13;
assign _c_doomhead[787] = 5'h13;
assign _c_doomhead[788] = 5'h13;
assign _c_doomhead[789] = 5'h0a;
assign _c_doomhead[790] = 5'h01;
assign _c_doomhead[791] = 5'h0e;
assign _c_doomhead[792] = 5'h00;
assign _c_doomhead[793] = 5'h00;
assign _c_doomhead[794] = 5'h00;
assign _c_doomhead[795] = 5'h00;
assign _c_doomhead[796] = 5'h00;
assign _c_doomhead[797] = 5'h00;
assign _c_doomhead[798] = 5'h00;
assign _c_doomhead[799] = 5'h00;
assign _c_doomhead[800] = 5'h00;
assign _c_doomhead[801] = 5'h00;
assign _c_doomhead[802] = 5'h00;
assign _c_doomhead[803] = 5'h00;
assign _c_doomhead[804] = 5'h00;
assign _c_doomhead[805] = 5'h00;
assign _c_doomhead[806] = 5'h00;
assign _c_doomhead[807] = 5'h04;
assign _c_doomhead[808] = 5'h0b;
assign _c_doomhead[809] = 5'h0c;
assign _c_doomhead[810] = 5'h14;
assign _c_doomhead[811] = 5'h13;
assign _c_doomhead[812] = 5'h0b;
assign _c_doomhead[813] = 5'h01;
assign _c_doomhead[814] = 5'h15;
assign _c_doomhead[815] = 5'h15;
assign _c_doomhead[816] = 5'h01;
assign _c_doomhead[817] = 5'h0b;
assign _c_doomhead[818] = 5'h13;
assign _c_doomhead[819] = 5'h14;
assign _c_doomhead[820] = 5'h0c;
assign _c_doomhead[821] = 5'h0b;
assign _c_doomhead[822] = 5'h04;
assign _c_doomhead[823] = 5'h00;
assign _c_doomhead[824] = 5'h00;
assign _c_doomhead[825] = 5'h00;
assign _c_doomhead[826] = 5'h00;
assign _c_doomhead[827] = 5'h00;
assign _c_doomhead[828] = 5'h00;
assign _c_doomhead[829] = 5'h00;
assign _c_doomhead[830] = 5'h00;
assign _c_doomhead[831] = 5'h00;
assign _c_doomhead[832] = 5'h00;
assign _c_doomhead[833] = 5'h00;
assign _c_doomhead[834] = 5'h00;
assign _c_doomhead[835] = 5'h00;
assign _c_doomhead[836] = 5'h00;
assign _c_doomhead[837] = 5'h00;
assign _c_doomhead[838] = 5'h00;
assign _c_doomhead[839] = 5'h00;
assign _c_doomhead[840] = 5'h04;
assign _c_doomhead[841] = 5'h0b;
assign _c_doomhead[842] = 5'h0c;
assign _c_doomhead[843] = 5'h14;
assign _c_doomhead[844] = 5'h13;
assign _c_doomhead[845] = 5'h13;
assign _c_doomhead[846] = 5'h12;
assign _c_doomhead[847] = 5'h12;
assign _c_doomhead[848] = 5'h13;
assign _c_doomhead[849] = 5'h13;
assign _c_doomhead[850] = 5'h14;
assign _c_doomhead[851] = 5'h0c;
assign _c_doomhead[852] = 5'h0b;
assign _c_doomhead[853] = 5'h04;
assign _c_doomhead[854] = 5'h00;
assign _c_doomhead[855] = 5'h00;
assign _c_doomhead[856] = 5'h00;
assign _c_doomhead[857] = 5'h00;
assign _c_doomhead[858] = 5'h00;
assign _c_doomhead[859] = 5'h00;
assign _c_doomhead[860] = 5'h00;
assign _c_doomhead[861] = 5'h00;
assign _c_doomhead[862] = 5'h00;
assign _c_doomhead[863] = 5'h00;
assign _c_doomhead[864] = 5'h00;
assign _c_doomhead[865] = 5'h00;
assign _c_doomhead[866] = 5'h00;
assign _c_doomhead[867] = 5'h00;
assign _c_doomhead[868] = 5'h00;
assign _c_doomhead[869] = 5'h00;
assign _c_doomhead[870] = 5'h00;
assign _c_doomhead[871] = 5'h00;
assign _c_doomhead[872] = 5'h00;
assign _c_doomhead[873] = 5'h0e;
assign _c_doomhead[874] = 5'h08;
assign _c_doomhead[875] = 5'h0a;
assign _c_doomhead[876] = 5'h0d;
assign _c_doomhead[877] = 5'h12;
assign _c_doomhead[878] = 5'h16;
assign _c_doomhead[879] = 5'h16;
assign _c_doomhead[880] = 5'h12;
assign _c_doomhead[881] = 5'h0d;
assign _c_doomhead[882] = 5'h0a;
assign _c_doomhead[883] = 5'h08;
assign _c_doomhead[884] = 5'h0e;
assign _c_doomhead[885] = 5'h00;
assign _c_doomhead[886] = 5'h00;
assign _c_doomhead[887] = 5'h00;
assign _c_doomhead[888] = 5'h00;
assign _c_doomhead[889] = 5'h00;
assign _c_doomhead[890] = 5'h00;
assign _c_doomhead[891] = 5'h00;
assign _c_doomhead[892] = 5'h00;
assign _c_doomhead[893] = 5'h00;
assign _c_doomhead[894] = 5'h00;
assign _c_doomhead[895] = 5'h00;
assign _c_doomhead[896] = 5'h00;
assign _c_doomhead[897] = 5'h00;
assign _c_doomhead[898] = 5'h00;
assign _c_doomhead[899] = 5'h00;
assign _c_doomhead[900] = 5'h00;
assign _c_doomhead[901] = 5'h00;
assign _c_doomhead[902] = 5'h00;
assign _c_doomhead[903] = 5'h00;
assign _c_doomhead[904] = 5'h00;
assign _c_doomhead[905] = 5'h00;
assign _c_doomhead[906] = 5'h00;
assign _c_doomhead[907] = 5'h04;
assign _c_doomhead[908] = 5'h01;
assign _c_doomhead[909] = 5'h09;
assign _c_doomhead[910] = 5'h09;
assign _c_doomhead[911] = 5'h09;
assign _c_doomhead[912] = 5'h09;
assign _c_doomhead[913] = 5'h01;
assign _c_doomhead[914] = 5'h04;
assign _c_doomhead[915] = 5'h00;
assign _c_doomhead[916] = 5'h00;
assign _c_doomhead[917] = 5'h00;
assign _c_doomhead[918] = 5'h00;
assign _c_doomhead[919] = 5'h00;
assign _c_doomhead[920] = 5'h00;
assign _c_doomhead[921] = 5'h00;
assign _c_doomhead[922] = 5'h00;
assign _c_doomhead[923] = 5'h00;
assign _c_doomhead[924] = 5'h00;
assign _c_doomhead[925] = 5'h00;
assign _c_doomhead[926] = 5'h00;
assign _c_doomhead[927] = 5'h00;
assign _c_doomhead[928] = 5'h00;
assign _c_doomhead[929] = 5'h00;
assign _c_doomhead[930] = 5'h00;
assign _c_doomhead[931] = 5'h00;
assign _c_doomhead[932] = 5'h00;
assign _c_doomhead[933] = 5'h00;
assign _c_doomhead[934] = 5'h00;
assign _c_doomhead[935] = 5'h00;
assign _c_doomhead[936] = 5'h00;
assign _c_doomhead[937] = 5'h00;
assign _c_doomhead[938] = 5'h00;
assign _c_doomhead[939] = 5'h00;
assign _c_doomhead[940] = 5'h00;
assign _c_doomhead[941] = 5'h00;
assign _c_doomhead[942] = 5'h00;
assign _c_doomhead[943] = 5'h00;
assign _c_doomhead[944] = 5'h00;
assign _c_doomhead[945] = 5'h00;
assign _c_doomhead[946] = 5'h00;
assign _c_doomhead[947] = 5'h00;
assign _c_doomhead[948] = 5'h00;
assign _c_doomhead[949] = 5'h00;
assign _c_doomhead[950] = 5'h00;
assign _c_doomhead[951] = 5'h00;
assign _c_doomhead[952] = 5'h00;
assign _c_doomhead[953] = 5'h00;
assign _c_doomhead[954] = 5'h00;
assign _c_doomhead[955] = 5'h00;
assign _c_doomhead[956] = 5'h00;
assign _c_doomhead[957] = 5'h00;
assign _c_doomhead[958] = 5'h00;
assign _c_doomhead[959] = 5'h00;
assign _c_doomhead[960] = 5'h00;
assign _c_doomhead[961] = 5'h00;
assign _c_doomhead[962] = 5'h00;
assign _c_doomhead[963] = 5'h00;
assign _c_doomhead[964] = 5'h00;
assign _c_doomhead[965] = 5'h00;
assign _c_doomhead[966] = 5'h00;
assign _c_doomhead[967] = 5'h00;
assign _c_doomhead[968] = 5'h00;
assign _c_doomhead[969] = 5'h00;
assign _c_doomhead[970] = 5'h00;
assign _c_doomhead[971] = 5'h00;
assign _c_doomhead[972] = 5'h00;
assign _c_doomhead[973] = 5'h00;
assign _c_doomhead[974] = 5'h00;
assign _c_doomhead[975] = 5'h00;
assign _c_doomhead[976] = 5'h00;
assign _c_doomhead[977] = 5'h00;
assign _c_doomhead[978] = 5'h00;
assign _c_doomhead[979] = 5'h00;
assign _c_doomhead[980] = 5'h00;
assign _c_doomhead[981] = 5'h00;
assign _c_doomhead[982] = 5'h00;
assign _c_doomhead[983] = 5'h00;
assign _c_doomhead[984] = 5'h00;
assign _c_doomhead[985] = 5'h00;
assign _c_doomhead[986] = 5'h00;
assign _c_doomhead[987] = 5'h00;
assign _c_doomhead[988] = 5'h00;
assign _c_doomhead[989] = 5'h00;
assign _c_doomhead[990] = 5'h00;
assign _c_doomhead[991] = 5'h00;
assign _c_doomhead[992] = 5'h00;
assign _c_doomhead[993] = 5'h00;
assign _c_doomhead[994] = 5'h00;
assign _c_doomhead[995] = 5'h00;
assign _c_doomhead[996] = 5'h00;
assign _c_doomhead[997] = 5'h00;
assign _c_doomhead[998] = 5'h00;
assign _c_doomhead[999] = 5'h00;
assign _c_doomhead[1000] = 5'h00;
assign _c_doomhead[1001] = 5'h00;
assign _c_doomhead[1002] = 5'h00;
assign _c_doomhead[1003] = 5'h00;
assign _c_doomhead[1004] = 5'h00;
assign _c_doomhead[1005] = 5'h00;
assign _c_doomhead[1006] = 5'h00;
assign _c_doomhead[1007] = 5'h00;
assign _c_doomhead[1008] = 5'h00;
assign _c_doomhead[1009] = 5'h00;
assign _c_doomhead[1010] = 5'h00;
assign _c_doomhead[1011] = 5'h00;
assign _c_doomhead[1012] = 5'h00;
assign _c_doomhead[1013] = 5'h00;
assign _c_doomhead[1014] = 5'h00;
assign _c_doomhead[1015] = 5'h00;
assign _c_doomhead[1016] = 5'h00;
assign _c_doomhead[1017] = 5'h00;
assign _c_doomhead[1018] = 5'h00;
assign _c_doomhead[1019] = 5'h00;
assign _c_doomhead[1020] = 5'h00;
assign _c_doomhead[1021] = 5'h00;
assign _c_doomhead[1022] = 5'h00;
assign _c_doomhead[1023] = 5'h00;
assign _c_doomhead[1024] = 5'h00;
assign _c_doomhead[1025] = 5'h00;
assign _c_doomhead[1026] = 5'h00;
assign _c_doomhead[1027] = 5'h00;
assign _c_doomhead[1028] = 5'h00;
assign _c_doomhead[1029] = 5'h00;
assign _c_doomhead[1030] = 5'h00;
assign _c_doomhead[1031] = 5'h00;
assign _c_doomhead[1032] = 5'h05;
assign _c_doomhead[1033] = 5'h02;
assign _c_doomhead[1034] = 5'h02;
assign _c_doomhead[1035] = 5'h02;
assign _c_doomhead[1036] = 5'h04;
assign _c_doomhead[1037] = 5'h06;
assign _c_doomhead[1038] = 5'h06;
assign _c_doomhead[1039] = 5'h06;
assign _c_doomhead[1040] = 5'h06;
assign _c_doomhead[1041] = 5'h06;
assign _c_doomhead[1042] = 5'h04;
assign _c_doomhead[1043] = 5'h02;
assign _c_doomhead[1044] = 5'h02;
assign _c_doomhead[1045] = 5'h05;
assign _c_doomhead[1046] = 5'h00;
assign _c_doomhead[1047] = 5'h00;
assign _c_doomhead[1048] = 5'h00;
assign _c_doomhead[1049] = 5'h00;
assign _c_doomhead[1050] = 5'h00;
assign _c_doomhead[1051] = 5'h00;
assign _c_doomhead[1052] = 5'h00;
assign _c_doomhead[1053] = 5'h00;
assign _c_doomhead[1054] = 5'h00;
assign _c_doomhead[1055] = 5'h00;
assign _c_doomhead[1056] = 5'h00;
assign _c_doomhead[1057] = 5'h00;
assign _c_doomhead[1058] = 5'h00;
assign _c_doomhead[1059] = 5'h00;
assign _c_doomhead[1060] = 5'h00;
assign _c_doomhead[1061] = 5'h00;
assign _c_doomhead[1062] = 5'h03;
assign _c_doomhead[1063] = 5'h02;
assign _c_doomhead[1064] = 5'h0e;
assign _c_doomhead[1065] = 5'h15;
assign _c_doomhead[1066] = 5'h01;
assign _c_doomhead[1067] = 5'h0b;
assign _c_doomhead[1068] = 5'h0f;
assign _c_doomhead[1069] = 5'h0c;
assign _c_doomhead[1070] = 5'h0c;
assign _c_doomhead[1071] = 5'h0c;
assign _c_doomhead[1072] = 5'h0f;
assign _c_doomhead[1073] = 5'h0b;
assign _c_doomhead[1074] = 5'h07;
assign _c_doomhead[1075] = 5'h06;
assign _c_doomhead[1076] = 5'h02;
assign _c_doomhead[1077] = 5'h0e;
assign _c_doomhead[1078] = 5'h02;
assign _c_doomhead[1079] = 5'h03;
assign _c_doomhead[1080] = 5'h00;
assign _c_doomhead[1081] = 5'h00;
assign _c_doomhead[1082] = 5'h00;
assign _c_doomhead[1083] = 5'h00;
assign _c_doomhead[1084] = 5'h00;
assign _c_doomhead[1085] = 5'h00;
assign _c_doomhead[1086] = 5'h00;
assign _c_doomhead[1087] = 5'h00;
assign _c_doomhead[1088] = 5'h00;
assign _c_doomhead[1089] = 5'h00;
assign _c_doomhead[1090] = 5'h00;
assign _c_doomhead[1091] = 5'h00;
assign _c_doomhead[1092] = 5'h00;
assign _c_doomhead[1093] = 5'h03;
assign _c_doomhead[1094] = 5'h02;
assign _c_doomhead[1095] = 5'h06;
assign _c_doomhead[1096] = 5'h01;
assign _c_doomhead[1097] = 5'h0b;
assign _c_doomhead[1098] = 5'h0f;
assign _c_doomhead[1099] = 5'h13;
assign _c_doomhead[1100] = 5'h0c;
assign _c_doomhead[1101] = 5'h0f;
assign _c_doomhead[1102] = 5'h0a;
assign _c_doomhead[1103] = 5'h07;
assign _c_doomhead[1104] = 5'h07;
assign _c_doomhead[1105] = 5'h07;
assign _c_doomhead[1106] = 5'h01;
assign _c_doomhead[1107] = 5'h01;
assign _c_doomhead[1108] = 5'h06;
assign _c_doomhead[1109] = 5'h06;
assign _c_doomhead[1110] = 5'h0e;
assign _c_doomhead[1111] = 5'h05;
assign _c_doomhead[1112] = 5'h03;
assign _c_doomhead[1113] = 5'h00;
assign _c_doomhead[1114] = 5'h00;
assign _c_doomhead[1115] = 5'h00;
assign _c_doomhead[1116] = 5'h00;
assign _c_doomhead[1117] = 5'h00;
assign _c_doomhead[1118] = 5'h00;
assign _c_doomhead[1119] = 5'h00;
assign _c_doomhead[1120] = 5'h00;
assign _c_doomhead[1121] = 5'h00;
assign _c_doomhead[1122] = 5'h00;
assign _c_doomhead[1123] = 5'h00;
assign _c_doomhead[1124] = 5'h00;
assign _c_doomhead[1125] = 5'h03;
assign _c_doomhead[1126] = 5'h06;
assign _c_doomhead[1127] = 5'h08;
assign _c_doomhead[1128] = 5'h06;
assign _c_doomhead[1129] = 5'h01;
assign _c_doomhead[1130] = 5'h07;
assign _c_doomhead[1131] = 5'h0a;
assign _c_doomhead[1132] = 5'h08;
assign _c_doomhead[1133] = 5'h0b;
assign _c_doomhead[1134] = 5'h01;
assign _c_doomhead[1135] = 5'h09;
assign _c_doomhead[1136] = 5'h06;
assign _c_doomhead[1137] = 5'h06;
assign _c_doomhead[1138] = 5'h06;
assign _c_doomhead[1139] = 5'h06;
assign _c_doomhead[1140] = 5'h02;
assign _c_doomhead[1141] = 5'h0e;
assign _c_doomhead[1142] = 5'h03;
assign _c_doomhead[1143] = 5'h03;
assign _c_doomhead[1144] = 5'h11;
assign _c_doomhead[1145] = 5'h00;
assign _c_doomhead[1146] = 5'h00;
assign _c_doomhead[1147] = 5'h00;
assign _c_doomhead[1148] = 5'h00;
assign _c_doomhead[1149] = 5'h00;
assign _c_doomhead[1150] = 5'h00;
assign _c_doomhead[1151] = 5'h00;
assign _c_doomhead[1152] = 5'h00;
assign _c_doomhead[1153] = 5'h00;
assign _c_doomhead[1154] = 5'h00;
assign _c_doomhead[1155] = 5'h00;
assign _c_doomhead[1156] = 5'h11;
assign _c_doomhead[1157] = 5'h10;
assign _c_doomhead[1158] = 5'h02;
assign _c_doomhead[1159] = 5'h06;
assign _c_doomhead[1160] = 5'h02;
assign _c_doomhead[1161] = 5'h01;
assign _c_doomhead[1162] = 5'h07;
assign _c_doomhead[1163] = 5'h01;
assign _c_doomhead[1164] = 5'h01;
assign _c_doomhead[1165] = 5'h01;
assign _c_doomhead[1166] = 5'h01;
assign _c_doomhead[1167] = 5'h05;
assign _c_doomhead[1168] = 5'h01;
assign _c_doomhead[1169] = 5'h02;
assign _c_doomhead[1170] = 5'h05;
assign _c_doomhead[1171] = 5'h02;
assign _c_doomhead[1172] = 5'h05;
assign _c_doomhead[1173] = 5'h03;
assign _c_doomhead[1174] = 5'h11;
assign _c_doomhead[1175] = 5'h11;
assign _c_doomhead[1176] = 5'h11;
assign _c_doomhead[1177] = 5'h11;
assign _c_doomhead[1178] = 5'h00;
assign _c_doomhead[1179] = 5'h00;
assign _c_doomhead[1180] = 5'h00;
assign _c_doomhead[1181] = 5'h00;
assign _c_doomhead[1182] = 5'h00;
assign _c_doomhead[1183] = 5'h00;
assign _c_doomhead[1184] = 5'h00;
assign _c_doomhead[1185] = 5'h00;
assign _c_doomhead[1186] = 5'h00;
assign _c_doomhead[1187] = 5'h00;
assign _c_doomhead[1188] = 5'h11;
assign _c_doomhead[1189] = 5'h10;
assign _c_doomhead[1190] = 5'h05;
assign _c_doomhead[1191] = 5'h0e;
assign _c_doomhead[1192] = 5'h02;
assign _c_doomhead[1193] = 5'h01;
assign _c_doomhead[1194] = 5'h0e;
assign _c_doomhead[1195] = 5'h07;
assign _c_doomhead[1196] = 5'h04;
assign _c_doomhead[1197] = 5'h04;
assign _c_doomhead[1198] = 5'h01;
assign _c_doomhead[1199] = 5'h04;
assign _c_doomhead[1200] = 5'h05;
assign _c_doomhead[1201] = 5'h04;
assign _c_doomhead[1202] = 5'h05;
assign _c_doomhead[1203] = 5'h10;
assign _c_doomhead[1204] = 5'h02;
assign _c_doomhead[1205] = 5'h11;
assign _c_doomhead[1206] = 5'h03;
assign _c_doomhead[1207] = 5'h03;
assign _c_doomhead[1208] = 5'h10;
assign _c_doomhead[1209] = 5'h11;
assign _c_doomhead[1210] = 5'h00;
assign _c_doomhead[1211] = 5'h00;
assign _c_doomhead[1212] = 5'h00;
assign _c_doomhead[1213] = 5'h00;
assign _c_doomhead[1214] = 5'h00;
assign _c_doomhead[1215] = 5'h00;
assign _c_doomhead[1216] = 5'h00;
assign _c_doomhead[1217] = 5'h00;
assign _c_doomhead[1218] = 5'h00;
assign _c_doomhead[1219] = 5'h00;
assign _c_doomhead[1220] = 5'h11;
assign _c_doomhead[1221] = 5'h05;
assign _c_doomhead[1222] = 5'h05;
assign _c_doomhead[1223] = 5'h06;
assign _c_doomhead[1224] = 5'h06;
assign _c_doomhead[1225] = 5'h0e;
assign _c_doomhead[1226] = 5'h01;
assign _c_doomhead[1227] = 5'h0e;
assign _c_doomhead[1228] = 5'h04;
assign _c_doomhead[1229] = 5'h06;
assign _c_doomhead[1230] = 5'h04;
assign _c_doomhead[1231] = 5'h04;
assign _c_doomhead[1232] = 5'h01;
assign _c_doomhead[1233] = 5'h01;
assign _c_doomhead[1234] = 5'h01;
assign _c_doomhead[1235] = 5'h08;
assign _c_doomhead[1236] = 5'h08;
assign _c_doomhead[1237] = 5'h04;
assign _c_doomhead[1238] = 5'h05;
assign _c_doomhead[1239] = 5'h10;
assign _c_doomhead[1240] = 5'h05;
assign _c_doomhead[1241] = 5'h11;
assign _c_doomhead[1242] = 5'h00;
assign _c_doomhead[1243] = 5'h00;
assign _c_doomhead[1244] = 5'h00;
assign _c_doomhead[1245] = 5'h00;
assign _c_doomhead[1246] = 5'h00;
assign _c_doomhead[1247] = 5'h00;
assign _c_doomhead[1248] = 5'h00;
assign _c_doomhead[1249] = 5'h00;
assign _c_doomhead[1250] = 5'h00;
assign _c_doomhead[1251] = 5'h00;
assign _c_doomhead[1252] = 5'h11;
assign _c_doomhead[1253] = 5'h05;
assign _c_doomhead[1254] = 5'h0e;
assign _c_doomhead[1255] = 5'h06;
assign _c_doomhead[1256] = 5'h01;
assign _c_doomhead[1257] = 5'h06;
assign _c_doomhead[1258] = 5'h0e;
assign _c_doomhead[1259] = 5'h09;
assign _c_doomhead[1260] = 5'h0e;
assign _c_doomhead[1261] = 5'h06;
assign _c_doomhead[1262] = 5'h01;
assign _c_doomhead[1263] = 5'h09;
assign _c_doomhead[1264] = 5'h0a;
assign _c_doomhead[1265] = 5'h07;
assign _c_doomhead[1266] = 5'h09;
assign _c_doomhead[1267] = 5'h01;
assign _c_doomhead[1268] = 5'h01;
assign _c_doomhead[1269] = 5'h01;
assign _c_doomhead[1270] = 5'h04;
assign _c_doomhead[1271] = 5'h05;
assign _c_doomhead[1272] = 5'h05;
assign _c_doomhead[1273] = 5'h11;
assign _c_doomhead[1274] = 5'h00;
assign _c_doomhead[1275] = 5'h00;
assign _c_doomhead[1276] = 5'h00;
assign _c_doomhead[1277] = 5'h00;
assign _c_doomhead[1278] = 5'h00;
assign _c_doomhead[1279] = 5'h00;
assign _c_doomhead[1280] = 5'h00;
assign _c_doomhead[1281] = 5'h00;
assign _c_doomhead[1282] = 5'h00;
assign _c_doomhead[1283] = 5'h00;
assign _c_doomhead[1284] = 5'h11;
assign _c_doomhead[1285] = 5'h05;
assign _c_doomhead[1286] = 5'h02;
assign _c_doomhead[1287] = 5'h01;
assign _c_doomhead[1288] = 5'h0b;
assign _c_doomhead[1289] = 5'h0a;
assign _c_doomhead[1290] = 5'h09;
assign _c_doomhead[1291] = 5'h09;
assign _c_doomhead[1292] = 5'h0a;
assign _c_doomhead[1293] = 5'h0a;
assign _c_doomhead[1294] = 5'h0a;
assign _c_doomhead[1295] = 5'h0a;
assign _c_doomhead[1296] = 5'h0a;
assign _c_doomhead[1297] = 5'h0a;
assign _c_doomhead[1298] = 5'h09;
assign _c_doomhead[1299] = 5'h09;
assign _c_doomhead[1300] = 5'h0a;
assign _c_doomhead[1301] = 5'h0b;
assign _c_doomhead[1302] = 5'h01;
assign _c_doomhead[1303] = 5'h0e;
assign _c_doomhead[1304] = 5'h05;
assign _c_doomhead[1305] = 5'h11;
assign _c_doomhead[1306] = 5'h00;
assign _c_doomhead[1307] = 5'h00;
assign _c_doomhead[1308] = 5'h00;
assign _c_doomhead[1309] = 5'h00;
assign _c_doomhead[1310] = 5'h00;
assign _c_doomhead[1311] = 5'h00;
assign _c_doomhead[1312] = 5'h00;
assign _c_doomhead[1313] = 5'h00;
assign _c_doomhead[1314] = 5'h00;
assign _c_doomhead[1315] = 5'h00;
assign _c_doomhead[1316] = 5'h11;
assign _c_doomhead[1317] = 5'h05;
assign _c_doomhead[1318] = 5'h06;
assign _c_doomhead[1319] = 5'h07;
assign _c_doomhead[1320] = 5'h0c;
assign _c_doomhead[1321] = 5'h13;
assign _c_doomhead[1322] = 5'h13;
assign _c_doomhead[1323] = 5'h0a;
assign _c_doomhead[1324] = 5'h09;
assign _c_doomhead[1325] = 5'h0b;
assign _c_doomhead[1326] = 5'h0b;
assign _c_doomhead[1327] = 5'h0b;
assign _c_doomhead[1328] = 5'h0b;
assign _c_doomhead[1329] = 5'h09;
assign _c_doomhead[1330] = 5'h0a;
assign _c_doomhead[1331] = 5'h13;
assign _c_doomhead[1332] = 5'h13;
assign _c_doomhead[1333] = 5'h0c;
assign _c_doomhead[1334] = 5'h07;
assign _c_doomhead[1335] = 5'h02;
assign _c_doomhead[1336] = 5'h05;
assign _c_doomhead[1337] = 5'h11;
assign _c_doomhead[1338] = 5'h00;
assign _c_doomhead[1339] = 5'h00;
assign _c_doomhead[1340] = 5'h00;
assign _c_doomhead[1341] = 5'h00;
assign _c_doomhead[1342] = 5'h00;
assign _c_doomhead[1343] = 5'h00;
assign _c_doomhead[1344] = 5'h00;
assign _c_doomhead[1345] = 5'h00;
assign _c_doomhead[1346] = 5'h00;
assign _c_doomhead[1347] = 5'h00;
assign _c_doomhead[1348] = 5'h11;
assign _c_doomhead[1349] = 5'h05;
assign _c_doomhead[1350] = 5'h06;
assign _c_doomhead[1351] = 5'h07;
assign _c_doomhead[1352] = 5'h0c;
assign _c_doomhead[1353] = 5'h19;
assign _c_doomhead[1354] = 5'h12;
assign _c_doomhead[1355] = 5'h0c;
assign _c_doomhead[1356] = 5'h0f;
assign _c_doomhead[1357] = 5'h09;
assign _c_doomhead[1358] = 5'h01;
assign _c_doomhead[1359] = 5'h01;
assign _c_doomhead[1360] = 5'h09;
assign _c_doomhead[1361] = 5'h0f;
assign _c_doomhead[1362] = 5'h0c;
assign _c_doomhead[1363] = 5'h12;
assign _c_doomhead[1364] = 5'h19;
assign _c_doomhead[1365] = 5'h0c;
assign _c_doomhead[1366] = 5'h07;
assign _c_doomhead[1367] = 5'h06;
assign _c_doomhead[1368] = 5'h05;
assign _c_doomhead[1369] = 5'h11;
assign _c_doomhead[1370] = 5'h00;
assign _c_doomhead[1371] = 5'h00;
assign _c_doomhead[1372] = 5'h00;
assign _c_doomhead[1373] = 5'h00;
assign _c_doomhead[1374] = 5'h00;
assign _c_doomhead[1375] = 5'h00;
assign _c_doomhead[1376] = 5'h00;
assign _c_doomhead[1377] = 5'h00;
assign _c_doomhead[1378] = 5'h00;
assign _c_doomhead[1379] = 5'h00;
assign _c_doomhead[1380] = 5'h11;
assign _c_doomhead[1381] = 5'h05;
assign _c_doomhead[1382] = 5'h06;
assign _c_doomhead[1383] = 5'h0a;
assign _c_doomhead[1384] = 5'h12;
assign _c_doomhead[1385] = 5'h16;
assign _c_doomhead[1386] = 5'h16;
assign _c_doomhead[1387] = 5'h12;
assign _c_doomhead[1388] = 5'h12;
assign _c_doomhead[1389] = 5'h0c;
assign _c_doomhead[1390] = 5'h0d;
assign _c_doomhead[1391] = 5'h0d;
assign _c_doomhead[1392] = 5'h0c;
assign _c_doomhead[1393] = 5'h12;
assign _c_doomhead[1394] = 5'h12;
assign _c_doomhead[1395] = 5'h07;
assign _c_doomhead[1396] = 5'h0e;
assign _c_doomhead[1397] = 5'h17;
assign _c_doomhead[1398] = 5'h10;
assign _c_doomhead[1399] = 5'h06;
assign _c_doomhead[1400] = 5'h05;
assign _c_doomhead[1401] = 5'h11;
assign _c_doomhead[1402] = 5'h00;
assign _c_doomhead[1403] = 5'h00;
assign _c_doomhead[1404] = 5'h00;
assign _c_doomhead[1405] = 5'h00;
assign _c_doomhead[1406] = 5'h00;
assign _c_doomhead[1407] = 5'h00;
assign _c_doomhead[1408] = 5'h00;
assign _c_doomhead[1409] = 5'h00;
assign _c_doomhead[1410] = 5'h00;
assign _c_doomhead[1411] = 5'h0a;
assign _c_doomhead[1412] = 5'h04;
assign _c_doomhead[1413] = 5'h05;
assign _c_doomhead[1414] = 5'h06;
assign _c_doomhead[1415] = 5'h10;
assign _c_doomhead[1416] = 5'h10;
assign _c_doomhead[1417] = 5'h0e;
assign _c_doomhead[1418] = 5'h09;
assign _c_doomhead[1419] = 5'h14;
assign _c_doomhead[1420] = 5'h16;
assign _c_doomhead[1421] = 5'h0f;
assign _c_doomhead[1422] = 5'h18;
assign _c_doomhead[1423] = 5'h18;
assign _c_doomhead[1424] = 5'h0f;
assign _c_doomhead[1425] = 5'h16;
assign _c_doomhead[1426] = 5'h07;
assign _c_doomhead[1427] = 5'h17;
assign _c_doomhead[1428] = 5'h10;
assign _c_doomhead[1429] = 5'h06;
assign _c_doomhead[1430] = 5'h08;
assign _c_doomhead[1431] = 5'h06;
assign _c_doomhead[1432] = 5'h05;
assign _c_doomhead[1433] = 5'h04;
assign _c_doomhead[1434] = 5'h0a;
assign _c_doomhead[1435] = 5'h00;
assign _c_doomhead[1436] = 5'h00;
assign _c_doomhead[1437] = 5'h00;
assign _c_doomhead[1438] = 5'h00;
assign _c_doomhead[1439] = 5'h00;
assign _c_doomhead[1440] = 5'h00;
assign _c_doomhead[1441] = 5'h00;
assign _c_doomhead[1442] = 5'h00;
assign _c_doomhead[1443] = 5'h0a;
assign _c_doomhead[1444] = 5'h04;
assign _c_doomhead[1445] = 5'h05;
assign _c_doomhead[1446] = 5'h0a;
assign _c_doomhead[1447] = 5'h08;
assign _c_doomhead[1448] = 5'h02;
assign _c_doomhead[1449] = 5'h10;
assign _c_doomhead[1450] = 5'h10;
assign _c_doomhead[1451] = 5'h10;
assign _c_doomhead[1452] = 5'h17;
assign _c_doomhead[1453] = 5'h02;
assign _c_doomhead[1454] = 5'h0b;
assign _c_doomhead[1455] = 5'h0b;
assign _c_doomhead[1456] = 5'h02;
assign _c_doomhead[1457] = 5'h17;
assign _c_doomhead[1458] = 5'h17;
assign _c_doomhead[1459] = 5'h17;
assign _c_doomhead[1460] = 5'h10;
assign _c_doomhead[1461] = 5'h02;
assign _c_doomhead[1462] = 5'h0a;
assign _c_doomhead[1463] = 5'h01;
assign _c_doomhead[1464] = 5'h05;
assign _c_doomhead[1465] = 5'h04;
assign _c_doomhead[1466] = 5'h0a;
assign _c_doomhead[1467] = 5'h00;
assign _c_doomhead[1468] = 5'h00;
assign _c_doomhead[1469] = 5'h00;
assign _c_doomhead[1470] = 5'h00;
assign _c_doomhead[1471] = 5'h00;
assign _c_doomhead[1472] = 5'h00;
assign _c_doomhead[1473] = 5'h00;
assign _c_doomhead[1474] = 5'h00;
assign _c_doomhead[1475] = 5'h01;
assign _c_doomhead[1476] = 5'h04;
assign _c_doomhead[1477] = 5'h04;
assign _c_doomhead[1478] = 5'h0a;
assign _c_doomhead[1479] = 5'h06;
assign _c_doomhead[1480] = 5'h00;
assign _c_doomhead[1481] = 5'h00;
assign _c_doomhead[1482] = 5'h07;
assign _c_doomhead[1483] = 5'h17;
assign _c_doomhead[1484] = 5'h17;
assign _c_doomhead[1485] = 5'h05;
assign _c_doomhead[1486] = 5'h0e;
assign _c_doomhead[1487] = 5'h0e;
assign _c_doomhead[1488] = 5'h05;
assign _c_doomhead[1489] = 5'h17;
assign _c_doomhead[1490] = 5'h15;
assign _c_doomhead[1491] = 5'h00;
assign _c_doomhead[1492] = 5'h07;
assign _c_doomhead[1493] = 5'h17;
assign _c_doomhead[1494] = 5'h06;
assign _c_doomhead[1495] = 5'h0a;
assign _c_doomhead[1496] = 5'h04;
assign _c_doomhead[1497] = 5'h04;
assign _c_doomhead[1498] = 5'h01;
assign _c_doomhead[1499] = 5'h00;
assign _c_doomhead[1500] = 5'h00;
assign _c_doomhead[1501] = 5'h00;
assign _c_doomhead[1502] = 5'h00;
assign _c_doomhead[1503] = 5'h00;
assign _c_doomhead[1504] = 5'h00;
assign _c_doomhead[1505] = 5'h00;
assign _c_doomhead[1506] = 5'h00;
assign _c_doomhead[1507] = 5'h04;
assign _c_doomhead[1508] = 5'h02;
assign _c_doomhead[1509] = 5'h08;
assign _c_doomhead[1510] = 5'h0a;
assign _c_doomhead[1511] = 5'h01;
assign _c_doomhead[1512] = 5'h0b;
assign _c_doomhead[1513] = 5'h19;
assign _c_doomhead[1514] = 5'h0b;
assign _c_doomhead[1515] = 5'h04;
assign _c_doomhead[1516] = 5'h02;
assign _c_doomhead[1517] = 5'h01;
assign _c_doomhead[1518] = 5'h0c;
assign _c_doomhead[1519] = 5'h0c;
assign _c_doomhead[1520] = 5'h01;
assign _c_doomhead[1521] = 5'h02;
assign _c_doomhead[1522] = 5'h04;
assign _c_doomhead[1523] = 5'h0b;
assign _c_doomhead[1524] = 5'h19;
assign _c_doomhead[1525] = 5'h0b;
assign _c_doomhead[1526] = 5'h01;
assign _c_doomhead[1527] = 5'h0a;
assign _c_doomhead[1528] = 5'h08;
assign _c_doomhead[1529] = 5'h02;
assign _c_doomhead[1530] = 5'h04;
assign _c_doomhead[1531] = 5'h00;
assign _c_doomhead[1532] = 5'h00;
assign _c_doomhead[1533] = 5'h00;
assign _c_doomhead[1534] = 5'h00;
assign _c_doomhead[1535] = 5'h00;
assign _c_doomhead[1536] = 5'h00;
assign _c_doomhead[1537] = 5'h00;
assign _c_doomhead[1538] = 5'h00;
assign _c_doomhead[1539] = 5'h08;
assign _c_doomhead[1540] = 5'h02;
assign _c_doomhead[1541] = 5'h08;
assign _c_doomhead[1542] = 5'h0d;
assign _c_doomhead[1543] = 5'h0d;
assign _c_doomhead[1544] = 5'h0f;
assign _c_doomhead[1545] = 5'h0b;
assign _c_doomhead[1546] = 5'h01;
assign _c_doomhead[1547] = 5'h0b;
assign _c_doomhead[1548] = 5'h0c;
assign _c_doomhead[1549] = 5'h0b;
assign _c_doomhead[1550] = 5'h18;
assign _c_doomhead[1551] = 5'h18;
assign _c_doomhead[1552] = 5'h0b;
assign _c_doomhead[1553] = 5'h0c;
assign _c_doomhead[1554] = 5'h0b;
assign _c_doomhead[1555] = 5'h01;
assign _c_doomhead[1556] = 5'h0b;
assign _c_doomhead[1557] = 5'h0f;
assign _c_doomhead[1558] = 5'h0d;
assign _c_doomhead[1559] = 5'h0d;
assign _c_doomhead[1560] = 5'h08;
assign _c_doomhead[1561] = 5'h02;
assign _c_doomhead[1562] = 5'h08;
assign _c_doomhead[1563] = 5'h00;
assign _c_doomhead[1564] = 5'h00;
assign _c_doomhead[1565] = 5'h00;
assign _c_doomhead[1566] = 5'h00;
assign _c_doomhead[1567] = 5'h00;
assign _c_doomhead[1568] = 5'h00;
assign _c_doomhead[1569] = 5'h00;
assign _c_doomhead[1570] = 5'h00;
assign _c_doomhead[1571] = 5'h01;
assign _c_doomhead[1572] = 5'h02;
assign _c_doomhead[1573] = 5'h01;
assign _c_doomhead[1574] = 5'h0c;
assign _c_doomhead[1575] = 5'h14;
assign _c_doomhead[1576] = 5'h19;
assign _c_doomhead[1577] = 5'h14;
assign _c_doomhead[1578] = 5'h13;
assign _c_doomhead[1579] = 5'h12;
assign _c_doomhead[1580] = 5'h16;
assign _c_doomhead[1581] = 5'h12;
assign _c_doomhead[1582] = 5'h16;
assign _c_doomhead[1583] = 5'h16;
assign _c_doomhead[1584] = 5'h12;
assign _c_doomhead[1585] = 5'h16;
assign _c_doomhead[1586] = 5'h12;
assign _c_doomhead[1587] = 5'h13;
assign _c_doomhead[1588] = 5'h14;
assign _c_doomhead[1589] = 5'h19;
assign _c_doomhead[1590] = 5'h14;
assign _c_doomhead[1591] = 5'h0c;
assign _c_doomhead[1592] = 5'h01;
assign _c_doomhead[1593] = 5'h02;
assign _c_doomhead[1594] = 5'h01;
assign _c_doomhead[1595] = 5'h00;
assign _c_doomhead[1596] = 5'h00;
assign _c_doomhead[1597] = 5'h00;
assign _c_doomhead[1598] = 5'h00;
assign _c_doomhead[1599] = 5'h00;
assign _c_doomhead[1600] = 5'h00;
assign _c_doomhead[1601] = 5'h00;
assign _c_doomhead[1602] = 5'h00;
assign _c_doomhead[1603] = 5'h00;
assign _c_doomhead[1604] = 5'h02;
assign _c_doomhead[1605] = 5'h08;
assign _c_doomhead[1606] = 5'h09;
assign _c_doomhead[1607] = 5'h0b;
assign _c_doomhead[1608] = 5'h0f;
assign _c_doomhead[1609] = 5'h0d;
assign _c_doomhead[1610] = 5'h19;
assign _c_doomhead[1611] = 5'h18;
assign _c_doomhead[1612] = 5'h14;
assign _c_doomhead[1613] = 5'h0d;
assign _c_doomhead[1614] = 5'h18;
assign _c_doomhead[1615] = 5'h16;
assign _c_doomhead[1616] = 5'h0d;
assign _c_doomhead[1617] = 5'h14;
assign _c_doomhead[1618] = 5'h18;
assign _c_doomhead[1619] = 5'h19;
assign _c_doomhead[1620] = 5'h0d;
assign _c_doomhead[1621] = 5'h0f;
assign _c_doomhead[1622] = 5'h0b;
assign _c_doomhead[1623] = 5'h09;
assign _c_doomhead[1624] = 5'h08;
assign _c_doomhead[1625] = 5'h02;
assign _c_doomhead[1626] = 5'h00;
assign _c_doomhead[1627] = 5'h00;
assign _c_doomhead[1628] = 5'h00;
assign _c_doomhead[1629] = 5'h00;
assign _c_doomhead[1630] = 5'h00;
assign _c_doomhead[1631] = 5'h00;
assign _c_doomhead[1632] = 5'h00;
assign _c_doomhead[1633] = 5'h00;
assign _c_doomhead[1634] = 5'h00;
assign _c_doomhead[1635] = 5'h00;
assign _c_doomhead[1636] = 5'h02;
assign _c_doomhead[1637] = 5'h06;
assign _c_doomhead[1638] = 5'h07;
assign _c_doomhead[1639] = 5'h09;
assign _c_doomhead[1640] = 5'h0f;
assign _c_doomhead[1641] = 5'h19;
assign _c_doomhead[1642] = 5'h16;
assign _c_doomhead[1643] = 5'h0d;
assign _c_doomhead[1644] = 5'h0b;
assign _c_doomhead[1645] = 5'h07;
assign _c_doomhead[1646] = 5'h00;
assign _c_doomhead[1647] = 5'h00;
assign _c_doomhead[1648] = 5'h07;
assign _c_doomhead[1649] = 5'h0b;
assign _c_doomhead[1650] = 5'h0d;
assign _c_doomhead[1651] = 5'h16;
assign _c_doomhead[1652] = 5'h19;
assign _c_doomhead[1653] = 5'h0f;
assign _c_doomhead[1654] = 5'h09;
assign _c_doomhead[1655] = 5'h07;
assign _c_doomhead[1656] = 5'h06;
assign _c_doomhead[1657] = 5'h02;
assign _c_doomhead[1658] = 5'h00;
assign _c_doomhead[1659] = 5'h00;
assign _c_doomhead[1660] = 5'h00;
assign _c_doomhead[1661] = 5'h00;
assign _c_doomhead[1662] = 5'h00;
assign _c_doomhead[1663] = 5'h00;
assign _c_doomhead[1664] = 5'h00;
assign _c_doomhead[1665] = 5'h00;
assign _c_doomhead[1666] = 5'h00;
assign _c_doomhead[1667] = 5'h00;
assign _c_doomhead[1668] = 5'h00;
assign _c_doomhead[1669] = 5'h06;
assign _c_doomhead[1670] = 5'h0a;
assign _c_doomhead[1671] = 5'h07;
assign _c_doomhead[1672] = 5'h0d;
assign _c_doomhead[1673] = 5'h16;
assign _c_doomhead[1674] = 5'h12;
assign _c_doomhead[1675] = 5'h09;
assign _c_doomhead[1676] = 5'h0e;
assign _c_doomhead[1677] = 5'h06;
assign _c_doomhead[1678] = 5'h08;
assign _c_doomhead[1679] = 5'h08;
assign _c_doomhead[1680] = 5'h06;
assign _c_doomhead[1681] = 5'h0e;
assign _c_doomhead[1682] = 5'h09;
assign _c_doomhead[1683] = 5'h12;
assign _c_doomhead[1684] = 5'h16;
assign _c_doomhead[1685] = 5'h0d;
assign _c_doomhead[1686] = 5'h07;
assign _c_doomhead[1687] = 5'h0a;
assign _c_doomhead[1688] = 5'h06;
assign _c_doomhead[1689] = 5'h00;
assign _c_doomhead[1690] = 5'h00;
assign _c_doomhead[1691] = 5'h00;
assign _c_doomhead[1692] = 5'h00;
assign _c_doomhead[1693] = 5'h00;
assign _c_doomhead[1694] = 5'h00;
assign _c_doomhead[1695] = 5'h00;
assign _c_doomhead[1696] = 5'h00;
assign _c_doomhead[1697] = 5'h00;
assign _c_doomhead[1698] = 5'h00;
assign _c_doomhead[1699] = 5'h00;
assign _c_doomhead[1700] = 5'h00;
assign _c_doomhead[1701] = 5'h02;
assign _c_doomhead[1702] = 5'h13;
assign _c_doomhead[1703] = 5'h07;
assign _c_doomhead[1704] = 5'h12;
assign _c_doomhead[1705] = 5'h18;
assign _c_doomhead[1706] = 5'h0f;
assign _c_doomhead[1707] = 5'h0c;
assign _c_doomhead[1708] = 5'h14;
assign _c_doomhead[1709] = 5'h0f;
assign _c_doomhead[1710] = 5'h09;
assign _c_doomhead[1711] = 5'h09;
assign _c_doomhead[1712] = 5'h0f;
assign _c_doomhead[1713] = 5'h14;
assign _c_doomhead[1714] = 5'h0c;
assign _c_doomhead[1715] = 5'h0f;
assign _c_doomhead[1716] = 5'h18;
assign _c_doomhead[1717] = 5'h12;
assign _c_doomhead[1718] = 5'h07;
assign _c_doomhead[1719] = 5'h13;
assign _c_doomhead[1720] = 5'h02;
assign _c_doomhead[1721] = 5'h00;
assign _c_doomhead[1722] = 5'h00;
assign _c_doomhead[1723] = 5'h00;
assign _c_doomhead[1724] = 5'h00;
assign _c_doomhead[1725] = 5'h00;
assign _c_doomhead[1726] = 5'h00;
assign _c_doomhead[1727] = 5'h00;
assign _c_doomhead[1728] = 5'h00;
assign _c_doomhead[1729] = 5'h00;
assign _c_doomhead[1730] = 5'h00;
assign _c_doomhead[1731] = 5'h00;
assign _c_doomhead[1732] = 5'h00;
assign _c_doomhead[1733] = 5'h0e;
assign _c_doomhead[1734] = 5'h0b;
assign _c_doomhead[1735] = 5'h09;
assign _c_doomhead[1736] = 5'h0d;
assign _c_doomhead[1737] = 5'h12;
assign _c_doomhead[1738] = 5'h0c;
assign _c_doomhead[1739] = 5'h0d;
assign _c_doomhead[1740] = 5'h18;
assign _c_doomhead[1741] = 5'h16;
assign _c_doomhead[1742] = 5'h0d;
assign _c_doomhead[1743] = 5'h0d;
assign _c_doomhead[1744] = 5'h16;
assign _c_doomhead[1745] = 5'h18;
assign _c_doomhead[1746] = 5'h0d;
assign _c_doomhead[1747] = 5'h0c;
assign _c_doomhead[1748] = 5'h12;
assign _c_doomhead[1749] = 5'h0d;
assign _c_doomhead[1750] = 5'h09;
assign _c_doomhead[1751] = 5'h0b;
assign _c_doomhead[1752] = 5'h0e;
assign _c_doomhead[1753] = 5'h00;
assign _c_doomhead[1754] = 5'h00;
assign _c_doomhead[1755] = 5'h00;
assign _c_doomhead[1756] = 5'h00;
assign _c_doomhead[1757] = 5'h00;
assign _c_doomhead[1758] = 5'h00;
assign _c_doomhead[1759] = 5'h00;
assign _c_doomhead[1760] = 5'h00;
assign _c_doomhead[1761] = 5'h00;
assign _c_doomhead[1762] = 5'h00;
assign _c_doomhead[1763] = 5'h00;
assign _c_doomhead[1764] = 5'h00;
assign _c_doomhead[1765] = 5'h00;
assign _c_doomhead[1766] = 5'h08;
assign _c_doomhead[1767] = 5'h0b;
assign _c_doomhead[1768] = 5'h13;
assign _c_doomhead[1769] = 5'h0d;
assign _c_doomhead[1770] = 5'h01;
assign _c_doomhead[1771] = 5'h06;
assign _c_doomhead[1772] = 5'h1f;
assign _c_doomhead[1773] = 5'h1f;
assign _c_doomhead[1774] = 5'h1f;
assign _c_doomhead[1775] = 5'h1f;
assign _c_doomhead[1776] = 5'h1f;
assign _c_doomhead[1777] = 5'h1f;
assign _c_doomhead[1778] = 5'h06;
assign _c_doomhead[1779] = 5'h01;
assign _c_doomhead[1780] = 5'h0d;
assign _c_doomhead[1781] = 5'h13;
assign _c_doomhead[1782] = 5'h0b;
assign _c_doomhead[1783] = 5'h08;
assign _c_doomhead[1784] = 5'h00;
assign _c_doomhead[1785] = 5'h00;
assign _c_doomhead[1786] = 5'h00;
assign _c_doomhead[1787] = 5'h00;
assign _c_doomhead[1788] = 5'h00;
assign _c_doomhead[1789] = 5'h00;
assign _c_doomhead[1790] = 5'h00;
assign _c_doomhead[1791] = 5'h00;
assign _c_doomhead[1792] = 5'h00;
assign _c_doomhead[1793] = 5'h00;
assign _c_doomhead[1794] = 5'h00;
assign _c_doomhead[1795] = 5'h00;
assign _c_doomhead[1796] = 5'h00;
assign _c_doomhead[1797] = 5'h00;
assign _c_doomhead[1798] = 5'h0e;
assign _c_doomhead[1799] = 5'h01;
assign _c_doomhead[1800] = 5'h0a;
assign _c_doomhead[1801] = 5'h13;
assign _c_doomhead[1802] = 5'h13;
assign _c_doomhead[1803] = 5'h13;
assign _c_doomhead[1804] = 5'h0d;
assign _c_doomhead[1805] = 5'h12;
assign _c_doomhead[1806] = 5'h12;
assign _c_doomhead[1807] = 5'h12;
assign _c_doomhead[1808] = 5'h12;
assign _c_doomhead[1809] = 5'h0d;
assign _c_doomhead[1810] = 5'h13;
assign _c_doomhead[1811] = 5'h13;
assign _c_doomhead[1812] = 5'h13;
assign _c_doomhead[1813] = 5'h0a;
assign _c_doomhead[1814] = 5'h01;
assign _c_doomhead[1815] = 5'h0e;
assign _c_doomhead[1816] = 5'h00;
assign _c_doomhead[1817] = 5'h00;
assign _c_doomhead[1818] = 5'h00;
assign _c_doomhead[1819] = 5'h00;
assign _c_doomhead[1820] = 5'h00;
assign _c_doomhead[1821] = 5'h00;
assign _c_doomhead[1822] = 5'h00;
assign _c_doomhead[1823] = 5'h00;
assign _c_doomhead[1824] = 5'h00;
assign _c_doomhead[1825] = 5'h00;
assign _c_doomhead[1826] = 5'h00;
assign _c_doomhead[1827] = 5'h00;
assign _c_doomhead[1828] = 5'h00;
assign _c_doomhead[1829] = 5'h00;
assign _c_doomhead[1830] = 5'h00;
assign _c_doomhead[1831] = 5'h04;
assign _c_doomhead[1832] = 5'h07;
assign _c_doomhead[1833] = 5'h0c;
assign _c_doomhead[1834] = 5'h14;
assign _c_doomhead[1835] = 5'h13;
assign _c_doomhead[1836] = 5'h0b;
assign _c_doomhead[1837] = 5'h01;
assign _c_doomhead[1838] = 5'h15;
assign _c_doomhead[1839] = 5'h15;
assign _c_doomhead[1840] = 5'h01;
assign _c_doomhead[1841] = 5'h0b;
assign _c_doomhead[1842] = 5'h13;
assign _c_doomhead[1843] = 5'h14;
assign _c_doomhead[1844] = 5'h0c;
assign _c_doomhead[1845] = 5'h07;
assign _c_doomhead[1846] = 5'h04;
assign _c_doomhead[1847] = 5'h00;
assign _c_doomhead[1848] = 5'h00;
assign _c_doomhead[1849] = 5'h00;
assign _c_doomhead[1850] = 5'h00;
assign _c_doomhead[1851] = 5'h00;
assign _c_doomhead[1852] = 5'h00;
assign _c_doomhead[1853] = 5'h00;
assign _c_doomhead[1854] = 5'h00;
assign _c_doomhead[1855] = 5'h00;
assign _c_doomhead[1856] = 5'h00;
assign _c_doomhead[1857] = 5'h00;
assign _c_doomhead[1858] = 5'h00;
assign _c_doomhead[1859] = 5'h00;
assign _c_doomhead[1860] = 5'h00;
assign _c_doomhead[1861] = 5'h00;
assign _c_doomhead[1862] = 5'h00;
assign _c_doomhead[1863] = 5'h00;
assign _c_doomhead[1864] = 5'h04;
assign _c_doomhead[1865] = 5'h09;
assign _c_doomhead[1866] = 5'h0c;
assign _c_doomhead[1867] = 5'h14;
assign _c_doomhead[1868] = 5'h13;
assign _c_doomhead[1869] = 5'h13;
assign _c_doomhead[1870] = 5'h12;
assign _c_doomhead[1871] = 5'h12;
assign _c_doomhead[1872] = 5'h13;
assign _c_doomhead[1873] = 5'h13;
assign _c_doomhead[1874] = 5'h14;
assign _c_doomhead[1875] = 5'h0c;
assign _c_doomhead[1876] = 5'h09;
assign _c_doomhead[1877] = 5'h04;
assign _c_doomhead[1878] = 5'h00;
assign _c_doomhead[1879] = 5'h00;
assign _c_doomhead[1880] = 5'h00;
assign _c_doomhead[1881] = 5'h00;
assign _c_doomhead[1882] = 5'h00;
assign _c_doomhead[1883] = 5'h00;
assign _c_doomhead[1884] = 5'h00;
assign _c_doomhead[1885] = 5'h00;
assign _c_doomhead[1886] = 5'h00;
assign _c_doomhead[1887] = 5'h00;
assign _c_doomhead[1888] = 5'h00;
assign _c_doomhead[1889] = 5'h00;
assign _c_doomhead[1890] = 5'h00;
assign _c_doomhead[1891] = 5'h00;
assign _c_doomhead[1892] = 5'h00;
assign _c_doomhead[1893] = 5'h00;
assign _c_doomhead[1894] = 5'h00;
assign _c_doomhead[1895] = 5'h00;
assign _c_doomhead[1896] = 5'h00;
assign _c_doomhead[1897] = 5'h0e;
assign _c_doomhead[1898] = 5'h08;
assign _c_doomhead[1899] = 5'h0a;
assign _c_doomhead[1900] = 5'h0d;
assign _c_doomhead[1901] = 5'h12;
assign _c_doomhead[1902] = 5'h16;
assign _c_doomhead[1903] = 5'h16;
assign _c_doomhead[1904] = 5'h12;
assign _c_doomhead[1905] = 5'h0d;
assign _c_doomhead[1906] = 5'h0a;
assign _c_doomhead[1907] = 5'h08;
assign _c_doomhead[1908] = 5'h0e;
assign _c_doomhead[1909] = 5'h00;
assign _c_doomhead[1910] = 5'h00;
assign _c_doomhead[1911] = 5'h00;
assign _c_doomhead[1912] = 5'h00;
assign _c_doomhead[1913] = 5'h00;
assign _c_doomhead[1914] = 5'h00;
assign _c_doomhead[1915] = 5'h00;
assign _c_doomhead[1916] = 5'h00;
assign _c_doomhead[1917] = 5'h00;
assign _c_doomhead[1918] = 5'h00;
assign _c_doomhead[1919] = 5'h00;
assign _c_doomhead[1920] = 5'h00;
assign _c_doomhead[1921] = 5'h00;
assign _c_doomhead[1922] = 5'h00;
assign _c_doomhead[1923] = 5'h00;
assign _c_doomhead[1924] = 5'h00;
assign _c_doomhead[1925] = 5'h00;
assign _c_doomhead[1926] = 5'h00;
assign _c_doomhead[1927] = 5'h00;
assign _c_doomhead[1928] = 5'h00;
assign _c_doomhead[1929] = 5'h00;
assign _c_doomhead[1930] = 5'h00;
assign _c_doomhead[1931] = 5'h04;
assign _c_doomhead[1932] = 5'h01;
assign _c_doomhead[1933] = 5'h09;
assign _c_doomhead[1934] = 5'h09;
assign _c_doomhead[1935] = 5'h09;
assign _c_doomhead[1936] = 5'h09;
assign _c_doomhead[1937] = 5'h01;
assign _c_doomhead[1938] = 5'h04;
assign _c_doomhead[1939] = 5'h00;
assign _c_doomhead[1940] = 5'h00;
assign _c_doomhead[1941] = 5'h00;
assign _c_doomhead[1942] = 5'h00;
assign _c_doomhead[1943] = 5'h00;
assign _c_doomhead[1944] = 5'h00;
assign _c_doomhead[1945] = 5'h00;
assign _c_doomhead[1946] = 5'h00;
assign _c_doomhead[1947] = 5'h00;
assign _c_doomhead[1948] = 5'h00;
assign _c_doomhead[1949] = 5'h00;
assign _c_doomhead[1950] = 5'h00;
assign _c_doomhead[1951] = 5'h00;
assign _c_doomhead[1952] = 5'h00;
assign _c_doomhead[1953] = 5'h00;
assign _c_doomhead[1954] = 5'h00;
assign _c_doomhead[1955] = 5'h00;
assign _c_doomhead[1956] = 5'h00;
assign _c_doomhead[1957] = 5'h00;
assign _c_doomhead[1958] = 5'h00;
assign _c_doomhead[1959] = 5'h00;
assign _c_doomhead[1960] = 5'h00;
assign _c_doomhead[1961] = 5'h00;
assign _c_doomhead[1962] = 5'h00;
assign _c_doomhead[1963] = 5'h00;
assign _c_doomhead[1964] = 5'h00;
assign _c_doomhead[1965] = 5'h00;
assign _c_doomhead[1966] = 5'h00;
assign _c_doomhead[1967] = 5'h00;
assign _c_doomhead[1968] = 5'h00;
assign _c_doomhead[1969] = 5'h00;
assign _c_doomhead[1970] = 5'h00;
assign _c_doomhead[1971] = 5'h00;
assign _c_doomhead[1972] = 5'h00;
assign _c_doomhead[1973] = 5'h00;
assign _c_doomhead[1974] = 5'h00;
assign _c_doomhead[1975] = 5'h00;
assign _c_doomhead[1976] = 5'h00;
assign _c_doomhead[1977] = 5'h00;
assign _c_doomhead[1978] = 5'h00;
assign _c_doomhead[1979] = 5'h00;
assign _c_doomhead[1980] = 5'h00;
assign _c_doomhead[1981] = 5'h00;
assign _c_doomhead[1982] = 5'h00;
assign _c_doomhead[1983] = 5'h00;
assign _c_doomhead[1984] = 5'h00;
assign _c_doomhead[1985] = 5'h00;
assign _c_doomhead[1986] = 5'h00;
assign _c_doomhead[1987] = 5'h00;
assign _c_doomhead[1988] = 5'h00;
assign _c_doomhead[1989] = 5'h00;
assign _c_doomhead[1990] = 5'h00;
assign _c_doomhead[1991] = 5'h00;
assign _c_doomhead[1992] = 5'h00;
assign _c_doomhead[1993] = 5'h00;
assign _c_doomhead[1994] = 5'h00;
assign _c_doomhead[1995] = 5'h00;
assign _c_doomhead[1996] = 5'h00;
assign _c_doomhead[1997] = 5'h00;
assign _c_doomhead[1998] = 5'h00;
assign _c_doomhead[1999] = 5'h00;
assign _c_doomhead[2000] = 5'h00;
assign _c_doomhead[2001] = 5'h00;
assign _c_doomhead[2002] = 5'h00;
assign _c_doomhead[2003] = 5'h00;
assign _c_doomhead[2004] = 5'h00;
assign _c_doomhead[2005] = 5'h00;
assign _c_doomhead[2006] = 5'h00;
assign _c_doomhead[2007] = 5'h00;
assign _c_doomhead[2008] = 5'h00;
assign _c_doomhead[2009] = 5'h00;
assign _c_doomhead[2010] = 5'h00;
assign _c_doomhead[2011] = 5'h00;
assign _c_doomhead[2012] = 5'h00;
assign _c_doomhead[2013] = 5'h00;
assign _c_doomhead[2014] = 5'h00;
assign _c_doomhead[2015] = 5'h00;
assign _c_doomhead[2016] = 5'h00;
assign _c_doomhead[2017] = 5'h00;
assign _c_doomhead[2018] = 5'h00;
assign _c_doomhead[2019] = 5'h00;
assign _c_doomhead[2020] = 5'h00;
assign _c_doomhead[2021] = 5'h00;
assign _c_doomhead[2022] = 5'h00;
assign _c_doomhead[2023] = 5'h00;
assign _c_doomhead[2024] = 5'h00;
assign _c_doomhead[2025] = 5'h00;
assign _c_doomhead[2026] = 5'h00;
assign _c_doomhead[2027] = 5'h00;
assign _c_doomhead[2028] = 5'h00;
assign _c_doomhead[2029] = 5'h00;
assign _c_doomhead[2030] = 5'h00;
assign _c_doomhead[2031] = 5'h00;
assign _c_doomhead[2032] = 5'h00;
assign _c_doomhead[2033] = 5'h00;
assign _c_doomhead[2034] = 5'h00;
assign _c_doomhead[2035] = 5'h00;
assign _c_doomhead[2036] = 5'h00;
assign _c_doomhead[2037] = 5'h00;
assign _c_doomhead[2038] = 5'h00;
assign _c_doomhead[2039] = 5'h00;
assign _c_doomhead[2040] = 5'h00;
assign _c_doomhead[2041] = 5'h00;
assign _c_doomhead[2042] = 5'h00;
assign _c_doomhead[2043] = 5'h00;
assign _c_doomhead[2044] = 5'h00;
assign _c_doomhead[2045] = 5'h00;
assign _c_doomhead[2046] = 5'h00;
assign _c_doomhead[2047] = 5'h00;
assign _c_doomhead[2048] = 5'h00;
assign _c_doomhead[2049] = 5'h00;
assign _c_doomhead[2050] = 5'h00;
assign _c_doomhead[2051] = 5'h00;
assign _c_doomhead[2052] = 5'h00;
assign _c_doomhead[2053] = 5'h00;
assign _c_doomhead[2054] = 5'h00;
assign _c_doomhead[2055] = 5'h00;
assign _c_doomhead[2056] = 5'h05;
assign _c_doomhead[2057] = 5'h02;
assign _c_doomhead[2058] = 5'h02;
assign _c_doomhead[2059] = 5'h02;
assign _c_doomhead[2060] = 5'h04;
assign _c_doomhead[2061] = 5'h06;
assign _c_doomhead[2062] = 5'h06;
assign _c_doomhead[2063] = 5'h06;
assign _c_doomhead[2064] = 5'h06;
assign _c_doomhead[2065] = 5'h06;
assign _c_doomhead[2066] = 5'h04;
assign _c_doomhead[2067] = 5'h02;
assign _c_doomhead[2068] = 5'h02;
assign _c_doomhead[2069] = 5'h05;
assign _c_doomhead[2070] = 5'h00;
assign _c_doomhead[2071] = 5'h00;
assign _c_doomhead[2072] = 5'h00;
assign _c_doomhead[2073] = 5'h00;
assign _c_doomhead[2074] = 5'h00;
assign _c_doomhead[2075] = 5'h00;
assign _c_doomhead[2076] = 5'h00;
assign _c_doomhead[2077] = 5'h00;
assign _c_doomhead[2078] = 5'h00;
assign _c_doomhead[2079] = 5'h00;
assign _c_doomhead[2080] = 5'h00;
assign _c_doomhead[2081] = 5'h00;
assign _c_doomhead[2082] = 5'h00;
assign _c_doomhead[2083] = 5'h00;
assign _c_doomhead[2084] = 5'h00;
assign _c_doomhead[2085] = 5'h00;
assign _c_doomhead[2086] = 5'h03;
assign _c_doomhead[2087] = 5'h02;
assign _c_doomhead[2088] = 5'h0e;
assign _c_doomhead[2089] = 5'h15;
assign _c_doomhead[2090] = 5'h01;
assign _c_doomhead[2091] = 5'h0b;
assign _c_doomhead[2092] = 5'h0f;
assign _c_doomhead[2093] = 5'h0c;
assign _c_doomhead[2094] = 5'h0c;
assign _c_doomhead[2095] = 5'h0c;
assign _c_doomhead[2096] = 5'h0f;
assign _c_doomhead[2097] = 5'h0b;
assign _c_doomhead[2098] = 5'h07;
assign _c_doomhead[2099] = 5'h06;
assign _c_doomhead[2100] = 5'h02;
assign _c_doomhead[2101] = 5'h0e;
assign _c_doomhead[2102] = 5'h02;
assign _c_doomhead[2103] = 5'h03;
assign _c_doomhead[2104] = 5'h00;
assign _c_doomhead[2105] = 5'h00;
assign _c_doomhead[2106] = 5'h00;
assign _c_doomhead[2107] = 5'h00;
assign _c_doomhead[2108] = 5'h00;
assign _c_doomhead[2109] = 5'h00;
assign _c_doomhead[2110] = 5'h00;
assign _c_doomhead[2111] = 5'h00;
assign _c_doomhead[2112] = 5'h00;
assign _c_doomhead[2113] = 5'h00;
assign _c_doomhead[2114] = 5'h00;
assign _c_doomhead[2115] = 5'h00;
assign _c_doomhead[2116] = 5'h00;
assign _c_doomhead[2117] = 5'h03;
assign _c_doomhead[2118] = 5'h02;
assign _c_doomhead[2119] = 5'h06;
assign _c_doomhead[2120] = 5'h01;
assign _c_doomhead[2121] = 5'h0b;
assign _c_doomhead[2122] = 5'h0f;
assign _c_doomhead[2123] = 5'h13;
assign _c_doomhead[2124] = 5'h0c;
assign _c_doomhead[2125] = 5'h0f;
assign _c_doomhead[2126] = 5'h0a;
assign _c_doomhead[2127] = 5'h07;
assign _c_doomhead[2128] = 5'h07;
assign _c_doomhead[2129] = 5'h07;
assign _c_doomhead[2130] = 5'h01;
assign _c_doomhead[2131] = 5'h01;
assign _c_doomhead[2132] = 5'h06;
assign _c_doomhead[2133] = 5'h06;
assign _c_doomhead[2134] = 5'h0e;
assign _c_doomhead[2135] = 5'h05;
assign _c_doomhead[2136] = 5'h03;
assign _c_doomhead[2137] = 5'h00;
assign _c_doomhead[2138] = 5'h00;
assign _c_doomhead[2139] = 5'h00;
assign _c_doomhead[2140] = 5'h00;
assign _c_doomhead[2141] = 5'h00;
assign _c_doomhead[2142] = 5'h00;
assign _c_doomhead[2143] = 5'h00;
assign _c_doomhead[2144] = 5'h00;
assign _c_doomhead[2145] = 5'h00;
assign _c_doomhead[2146] = 5'h00;
assign _c_doomhead[2147] = 5'h00;
assign _c_doomhead[2148] = 5'h00;
assign _c_doomhead[2149] = 5'h03;
assign _c_doomhead[2150] = 5'h06;
assign _c_doomhead[2151] = 5'h08;
assign _c_doomhead[2152] = 5'h06;
assign _c_doomhead[2153] = 5'h01;
assign _c_doomhead[2154] = 5'h07;
assign _c_doomhead[2155] = 5'h0a;
assign _c_doomhead[2156] = 5'h08;
assign _c_doomhead[2157] = 5'h0b;
assign _c_doomhead[2158] = 5'h01;
assign _c_doomhead[2159] = 5'h09;
assign _c_doomhead[2160] = 5'h06;
assign _c_doomhead[2161] = 5'h06;
assign _c_doomhead[2162] = 5'h06;
assign _c_doomhead[2163] = 5'h06;
assign _c_doomhead[2164] = 5'h02;
assign _c_doomhead[2165] = 5'h0e;
assign _c_doomhead[2166] = 5'h03;
assign _c_doomhead[2167] = 5'h03;
assign _c_doomhead[2168] = 5'h11;
assign _c_doomhead[2169] = 5'h00;
assign _c_doomhead[2170] = 5'h00;
assign _c_doomhead[2171] = 5'h00;
assign _c_doomhead[2172] = 5'h00;
assign _c_doomhead[2173] = 5'h00;
assign _c_doomhead[2174] = 5'h00;
assign _c_doomhead[2175] = 5'h00;
assign _c_doomhead[2176] = 5'h00;
assign _c_doomhead[2177] = 5'h00;
assign _c_doomhead[2178] = 5'h00;
assign _c_doomhead[2179] = 5'h00;
assign _c_doomhead[2180] = 5'h11;
assign _c_doomhead[2181] = 5'h10;
assign _c_doomhead[2182] = 5'h02;
assign _c_doomhead[2183] = 5'h06;
assign _c_doomhead[2184] = 5'h02;
assign _c_doomhead[2185] = 5'h01;
assign _c_doomhead[2186] = 5'h07;
assign _c_doomhead[2187] = 5'h01;
assign _c_doomhead[2188] = 5'h01;
assign _c_doomhead[2189] = 5'h01;
assign _c_doomhead[2190] = 5'h01;
assign _c_doomhead[2191] = 5'h05;
assign _c_doomhead[2192] = 5'h01;
assign _c_doomhead[2193] = 5'h02;
assign _c_doomhead[2194] = 5'h05;
assign _c_doomhead[2195] = 5'h02;
assign _c_doomhead[2196] = 5'h05;
assign _c_doomhead[2197] = 5'h03;
assign _c_doomhead[2198] = 5'h11;
assign _c_doomhead[2199] = 5'h11;
assign _c_doomhead[2200] = 5'h11;
assign _c_doomhead[2201] = 5'h11;
assign _c_doomhead[2202] = 5'h00;
assign _c_doomhead[2203] = 5'h00;
assign _c_doomhead[2204] = 5'h00;
assign _c_doomhead[2205] = 5'h00;
assign _c_doomhead[2206] = 5'h00;
assign _c_doomhead[2207] = 5'h00;
assign _c_doomhead[2208] = 5'h00;
assign _c_doomhead[2209] = 5'h00;
assign _c_doomhead[2210] = 5'h00;
assign _c_doomhead[2211] = 5'h00;
assign _c_doomhead[2212] = 5'h11;
assign _c_doomhead[2213] = 5'h10;
assign _c_doomhead[2214] = 5'h05;
assign _c_doomhead[2215] = 5'h0e;
assign _c_doomhead[2216] = 5'h02;
assign _c_doomhead[2217] = 5'h01;
assign _c_doomhead[2218] = 5'h0e;
assign _c_doomhead[2219] = 5'h07;
assign _c_doomhead[2220] = 5'h04;
assign _c_doomhead[2221] = 5'h04;
assign _c_doomhead[2222] = 5'h01;
assign _c_doomhead[2223] = 5'h04;
assign _c_doomhead[2224] = 5'h05;
assign _c_doomhead[2225] = 5'h04;
assign _c_doomhead[2226] = 5'h05;
assign _c_doomhead[2227] = 5'h10;
assign _c_doomhead[2228] = 5'h02;
assign _c_doomhead[2229] = 5'h11;
assign _c_doomhead[2230] = 5'h03;
assign _c_doomhead[2231] = 5'h03;
assign _c_doomhead[2232] = 5'h10;
assign _c_doomhead[2233] = 5'h11;
assign _c_doomhead[2234] = 5'h00;
assign _c_doomhead[2235] = 5'h00;
assign _c_doomhead[2236] = 5'h00;
assign _c_doomhead[2237] = 5'h00;
assign _c_doomhead[2238] = 5'h00;
assign _c_doomhead[2239] = 5'h00;
assign _c_doomhead[2240] = 5'h00;
assign _c_doomhead[2241] = 5'h00;
assign _c_doomhead[2242] = 5'h00;
assign _c_doomhead[2243] = 5'h00;
assign _c_doomhead[2244] = 5'h11;
assign _c_doomhead[2245] = 5'h05;
assign _c_doomhead[2246] = 5'h05;
assign _c_doomhead[2247] = 5'h06;
assign _c_doomhead[2248] = 5'h06;
assign _c_doomhead[2249] = 5'h0e;
assign _c_doomhead[2250] = 5'h01;
assign _c_doomhead[2251] = 5'h0e;
assign _c_doomhead[2252] = 5'h04;
assign _c_doomhead[2253] = 5'h06;
assign _c_doomhead[2254] = 5'h04;
assign _c_doomhead[2255] = 5'h04;
assign _c_doomhead[2256] = 5'h01;
assign _c_doomhead[2257] = 5'h01;
assign _c_doomhead[2258] = 5'h01;
assign _c_doomhead[2259] = 5'h08;
assign _c_doomhead[2260] = 5'h08;
assign _c_doomhead[2261] = 5'h04;
assign _c_doomhead[2262] = 5'h05;
assign _c_doomhead[2263] = 5'h10;
assign _c_doomhead[2264] = 5'h05;
assign _c_doomhead[2265] = 5'h11;
assign _c_doomhead[2266] = 5'h00;
assign _c_doomhead[2267] = 5'h00;
assign _c_doomhead[2268] = 5'h00;
assign _c_doomhead[2269] = 5'h00;
assign _c_doomhead[2270] = 5'h00;
assign _c_doomhead[2271] = 5'h00;
assign _c_doomhead[2272] = 5'h00;
assign _c_doomhead[2273] = 5'h00;
assign _c_doomhead[2274] = 5'h00;
assign _c_doomhead[2275] = 5'h00;
assign _c_doomhead[2276] = 5'h11;
assign _c_doomhead[2277] = 5'h05;
assign _c_doomhead[2278] = 5'h0e;
assign _c_doomhead[2279] = 5'h06;
assign _c_doomhead[2280] = 5'h01;
assign _c_doomhead[2281] = 5'h06;
assign _c_doomhead[2282] = 5'h0e;
assign _c_doomhead[2283] = 5'h09;
assign _c_doomhead[2284] = 5'h0e;
assign _c_doomhead[2285] = 5'h06;
assign _c_doomhead[2286] = 5'h01;
assign _c_doomhead[2287] = 5'h09;
assign _c_doomhead[2288] = 5'h0a;
assign _c_doomhead[2289] = 5'h07;
assign _c_doomhead[2290] = 5'h09;
assign _c_doomhead[2291] = 5'h01;
assign _c_doomhead[2292] = 5'h01;
assign _c_doomhead[2293] = 5'h01;
assign _c_doomhead[2294] = 5'h04;
assign _c_doomhead[2295] = 5'h05;
assign _c_doomhead[2296] = 5'h05;
assign _c_doomhead[2297] = 5'h11;
assign _c_doomhead[2298] = 5'h00;
assign _c_doomhead[2299] = 5'h00;
assign _c_doomhead[2300] = 5'h00;
assign _c_doomhead[2301] = 5'h00;
assign _c_doomhead[2302] = 5'h00;
assign _c_doomhead[2303] = 5'h00;
assign _c_doomhead[2304] = 5'h00;
assign _c_doomhead[2305] = 5'h00;
assign _c_doomhead[2306] = 5'h00;
assign _c_doomhead[2307] = 5'h00;
assign _c_doomhead[2308] = 5'h11;
assign _c_doomhead[2309] = 5'h05;
assign _c_doomhead[2310] = 5'h02;
assign _c_doomhead[2311] = 5'h01;
assign _c_doomhead[2312] = 5'h0b;
assign _c_doomhead[2313] = 5'h0a;
assign _c_doomhead[2314] = 5'h09;
assign _c_doomhead[2315] = 5'h09;
assign _c_doomhead[2316] = 5'h0a;
assign _c_doomhead[2317] = 5'h0a;
assign _c_doomhead[2318] = 5'h0a;
assign _c_doomhead[2319] = 5'h0a;
assign _c_doomhead[2320] = 5'h0a;
assign _c_doomhead[2321] = 5'h0a;
assign _c_doomhead[2322] = 5'h09;
assign _c_doomhead[2323] = 5'h09;
assign _c_doomhead[2324] = 5'h0a;
assign _c_doomhead[2325] = 5'h0b;
assign _c_doomhead[2326] = 5'h01;
assign _c_doomhead[2327] = 5'h0e;
assign _c_doomhead[2328] = 5'h05;
assign _c_doomhead[2329] = 5'h11;
assign _c_doomhead[2330] = 5'h00;
assign _c_doomhead[2331] = 5'h00;
assign _c_doomhead[2332] = 5'h00;
assign _c_doomhead[2333] = 5'h00;
assign _c_doomhead[2334] = 5'h00;
assign _c_doomhead[2335] = 5'h00;
assign _c_doomhead[2336] = 5'h00;
assign _c_doomhead[2337] = 5'h00;
assign _c_doomhead[2338] = 5'h00;
assign _c_doomhead[2339] = 5'h00;
assign _c_doomhead[2340] = 5'h11;
assign _c_doomhead[2341] = 5'h05;
assign _c_doomhead[2342] = 5'h06;
assign _c_doomhead[2343] = 5'h07;
assign _c_doomhead[2344] = 5'h0c;
assign _c_doomhead[2345] = 5'h13;
assign _c_doomhead[2346] = 5'h13;
assign _c_doomhead[2347] = 5'h0a;
assign _c_doomhead[2348] = 5'h09;
assign _c_doomhead[2349] = 5'h0b;
assign _c_doomhead[2350] = 5'h0b;
assign _c_doomhead[2351] = 5'h0b;
assign _c_doomhead[2352] = 5'h0b;
assign _c_doomhead[2353] = 5'h09;
assign _c_doomhead[2354] = 5'h0a;
assign _c_doomhead[2355] = 5'h13;
assign _c_doomhead[2356] = 5'h13;
assign _c_doomhead[2357] = 5'h0c;
assign _c_doomhead[2358] = 5'h07;
assign _c_doomhead[2359] = 5'h02;
assign _c_doomhead[2360] = 5'h05;
assign _c_doomhead[2361] = 5'h11;
assign _c_doomhead[2362] = 5'h00;
assign _c_doomhead[2363] = 5'h00;
assign _c_doomhead[2364] = 5'h00;
assign _c_doomhead[2365] = 5'h00;
assign _c_doomhead[2366] = 5'h00;
assign _c_doomhead[2367] = 5'h00;
assign _c_doomhead[2368] = 5'h00;
assign _c_doomhead[2369] = 5'h00;
assign _c_doomhead[2370] = 5'h00;
assign _c_doomhead[2371] = 5'h00;
assign _c_doomhead[2372] = 5'h11;
assign _c_doomhead[2373] = 5'h05;
assign _c_doomhead[2374] = 5'h06;
assign _c_doomhead[2375] = 5'h07;
assign _c_doomhead[2376] = 5'h0c;
assign _c_doomhead[2377] = 5'h19;
assign _c_doomhead[2378] = 5'h12;
assign _c_doomhead[2379] = 5'h0c;
assign _c_doomhead[2380] = 5'h0f;
assign _c_doomhead[2381] = 5'h09;
assign _c_doomhead[2382] = 5'h01;
assign _c_doomhead[2383] = 5'h01;
assign _c_doomhead[2384] = 5'h09;
assign _c_doomhead[2385] = 5'h0f;
assign _c_doomhead[2386] = 5'h0c;
assign _c_doomhead[2387] = 5'h12;
assign _c_doomhead[2388] = 5'h19;
assign _c_doomhead[2389] = 5'h0c;
assign _c_doomhead[2390] = 5'h07;
assign _c_doomhead[2391] = 5'h06;
assign _c_doomhead[2392] = 5'h05;
assign _c_doomhead[2393] = 5'h11;
assign _c_doomhead[2394] = 5'h00;
assign _c_doomhead[2395] = 5'h00;
assign _c_doomhead[2396] = 5'h00;
assign _c_doomhead[2397] = 5'h00;
assign _c_doomhead[2398] = 5'h00;
assign _c_doomhead[2399] = 5'h00;
assign _c_doomhead[2400] = 5'h00;
assign _c_doomhead[2401] = 5'h00;
assign _c_doomhead[2402] = 5'h00;
assign _c_doomhead[2403] = 5'h00;
assign _c_doomhead[2404] = 5'h11;
assign _c_doomhead[2405] = 5'h05;
assign _c_doomhead[2406] = 5'h06;
assign _c_doomhead[2407] = 5'h10;
assign _c_doomhead[2408] = 5'h17;
assign _c_doomhead[2409] = 5'h0e;
assign _c_doomhead[2410] = 5'h07;
assign _c_doomhead[2411] = 5'h12;
assign _c_doomhead[2412] = 5'h12;
assign _c_doomhead[2413] = 5'h0c;
assign _c_doomhead[2414] = 5'h0d;
assign _c_doomhead[2415] = 5'h0d;
assign _c_doomhead[2416] = 5'h0c;
assign _c_doomhead[2417] = 5'h12;
assign _c_doomhead[2418] = 5'h12;
assign _c_doomhead[2419] = 5'h16;
assign _c_doomhead[2420] = 5'h16;
assign _c_doomhead[2421] = 5'h12;
assign _c_doomhead[2422] = 5'h0a;
assign _c_doomhead[2423] = 5'h06;
assign _c_doomhead[2424] = 5'h05;
assign _c_doomhead[2425] = 5'h11;
assign _c_doomhead[2426] = 5'h00;
assign _c_doomhead[2427] = 5'h00;
assign _c_doomhead[2428] = 5'h00;
assign _c_doomhead[2429] = 5'h00;
assign _c_doomhead[2430] = 5'h00;
assign _c_doomhead[2431] = 5'h00;
assign _c_doomhead[2432] = 5'h00;
assign _c_doomhead[2433] = 5'h00;
assign _c_doomhead[2434] = 5'h00;
assign _c_doomhead[2435] = 5'h0a;
assign _c_doomhead[2436] = 5'h04;
assign _c_doomhead[2437] = 5'h05;
assign _c_doomhead[2438] = 5'h06;
assign _c_doomhead[2439] = 5'h08;
assign _c_doomhead[2440] = 5'h06;
assign _c_doomhead[2441] = 5'h10;
assign _c_doomhead[2442] = 5'h17;
assign _c_doomhead[2443] = 5'h07;
assign _c_doomhead[2444] = 5'h16;
assign _c_doomhead[2445] = 5'h0f;
assign _c_doomhead[2446] = 5'h18;
assign _c_doomhead[2447] = 5'h18;
assign _c_doomhead[2448] = 5'h0f;
assign _c_doomhead[2449] = 5'h16;
assign _c_doomhead[2450] = 5'h14;
assign _c_doomhead[2451] = 5'h09;
assign _c_doomhead[2452] = 5'h0e;
assign _c_doomhead[2453] = 5'h10;
assign _c_doomhead[2454] = 5'h10;
assign _c_doomhead[2455] = 5'h06;
assign _c_doomhead[2456] = 5'h05;
assign _c_doomhead[2457] = 5'h04;
assign _c_doomhead[2458] = 5'h0a;
assign _c_doomhead[2459] = 5'h00;
assign _c_doomhead[2460] = 5'h00;
assign _c_doomhead[2461] = 5'h00;
assign _c_doomhead[2462] = 5'h00;
assign _c_doomhead[2463] = 5'h00;
assign _c_doomhead[2464] = 5'h00;
assign _c_doomhead[2465] = 5'h00;
assign _c_doomhead[2466] = 5'h00;
assign _c_doomhead[2467] = 5'h0a;
assign _c_doomhead[2468] = 5'h04;
assign _c_doomhead[2469] = 5'h05;
assign _c_doomhead[2470] = 5'h01;
assign _c_doomhead[2471] = 5'h0a;
assign _c_doomhead[2472] = 5'h02;
assign _c_doomhead[2473] = 5'h10;
assign _c_doomhead[2474] = 5'h17;
assign _c_doomhead[2475] = 5'h17;
assign _c_doomhead[2476] = 5'h17;
assign _c_doomhead[2477] = 5'h02;
assign _c_doomhead[2478] = 5'h0b;
assign _c_doomhead[2479] = 5'h0b;
assign _c_doomhead[2480] = 5'h02;
assign _c_doomhead[2481] = 5'h17;
assign _c_doomhead[2482] = 5'h10;
assign _c_doomhead[2483] = 5'h10;
assign _c_doomhead[2484] = 5'h10;
assign _c_doomhead[2485] = 5'h02;
assign _c_doomhead[2486] = 5'h08;
assign _c_doomhead[2487] = 5'h0a;
assign _c_doomhead[2488] = 5'h05;
assign _c_doomhead[2489] = 5'h04;
assign _c_doomhead[2490] = 5'h0a;
assign _c_doomhead[2491] = 5'h00;
assign _c_doomhead[2492] = 5'h00;
assign _c_doomhead[2493] = 5'h00;
assign _c_doomhead[2494] = 5'h00;
assign _c_doomhead[2495] = 5'h00;
assign _c_doomhead[2496] = 5'h00;
assign _c_doomhead[2497] = 5'h00;
assign _c_doomhead[2498] = 5'h00;
assign _c_doomhead[2499] = 5'h01;
assign _c_doomhead[2500] = 5'h04;
assign _c_doomhead[2501] = 5'h04;
assign _c_doomhead[2502] = 5'h0a;
assign _c_doomhead[2503] = 5'h06;
assign _c_doomhead[2504] = 5'h17;
assign _c_doomhead[2505] = 5'h17;
assign _c_doomhead[2506] = 5'h00;
assign _c_doomhead[2507] = 5'h15;
assign _c_doomhead[2508] = 5'h17;
assign _c_doomhead[2509] = 5'h05;
assign _c_doomhead[2510] = 5'h0e;
assign _c_doomhead[2511] = 5'h0e;
assign _c_doomhead[2512] = 5'h05;
assign _c_doomhead[2513] = 5'h17;
assign _c_doomhead[2514] = 5'h17;
assign _c_doomhead[2515] = 5'h17;
assign _c_doomhead[2516] = 5'h00;
assign _c_doomhead[2517] = 5'h00;
assign _c_doomhead[2518] = 5'h06;
assign _c_doomhead[2519] = 5'h0a;
assign _c_doomhead[2520] = 5'h04;
assign _c_doomhead[2521] = 5'h04;
assign _c_doomhead[2522] = 5'h01;
assign _c_doomhead[2523] = 5'h00;
assign _c_doomhead[2524] = 5'h00;
assign _c_doomhead[2525] = 5'h00;
assign _c_doomhead[2526] = 5'h00;
assign _c_doomhead[2527] = 5'h00;
assign _c_doomhead[2528] = 5'h00;
assign _c_doomhead[2529] = 5'h00;
assign _c_doomhead[2530] = 5'h00;
assign _c_doomhead[2531] = 5'h04;
assign _c_doomhead[2532] = 5'h02;
assign _c_doomhead[2533] = 5'h08;
assign _c_doomhead[2534] = 5'h0a;
assign _c_doomhead[2535] = 5'h01;
assign _c_doomhead[2536] = 5'h0b;
assign _c_doomhead[2537] = 5'h19;
assign _c_doomhead[2538] = 5'h0b;
assign _c_doomhead[2539] = 5'h04;
assign _c_doomhead[2540] = 5'h02;
assign _c_doomhead[2541] = 5'h01;
assign _c_doomhead[2542] = 5'h0c;
assign _c_doomhead[2543] = 5'h0c;
assign _c_doomhead[2544] = 5'h01;
assign _c_doomhead[2545] = 5'h02;
assign _c_doomhead[2546] = 5'h04;
assign _c_doomhead[2547] = 5'h0b;
assign _c_doomhead[2548] = 5'h19;
assign _c_doomhead[2549] = 5'h0b;
assign _c_doomhead[2550] = 5'h01;
assign _c_doomhead[2551] = 5'h0a;
assign _c_doomhead[2552] = 5'h08;
assign _c_doomhead[2553] = 5'h02;
assign _c_doomhead[2554] = 5'h04;
assign _c_doomhead[2555] = 5'h00;
assign _c_doomhead[2556] = 5'h00;
assign _c_doomhead[2557] = 5'h00;
assign _c_doomhead[2558] = 5'h00;
assign _c_doomhead[2559] = 5'h00;
assign _c_doomhead[2560] = 5'h00;
assign _c_doomhead[2561] = 5'h00;
assign _c_doomhead[2562] = 5'h00;
assign _c_doomhead[2563] = 5'h08;
assign _c_doomhead[2564] = 5'h02;
assign _c_doomhead[2565] = 5'h08;
assign _c_doomhead[2566] = 5'h0d;
assign _c_doomhead[2567] = 5'h0d;
assign _c_doomhead[2568] = 5'h0f;
assign _c_doomhead[2569] = 5'h0b;
assign _c_doomhead[2570] = 5'h01;
assign _c_doomhead[2571] = 5'h0b;
assign _c_doomhead[2572] = 5'h0c;
assign _c_doomhead[2573] = 5'h0b;
assign _c_doomhead[2574] = 5'h18;
assign _c_doomhead[2575] = 5'h18;
assign _c_doomhead[2576] = 5'h0b;
assign _c_doomhead[2577] = 5'h0c;
assign _c_doomhead[2578] = 5'h0b;
assign _c_doomhead[2579] = 5'h01;
assign _c_doomhead[2580] = 5'h0b;
assign _c_doomhead[2581] = 5'h0f;
assign _c_doomhead[2582] = 5'h0d;
assign _c_doomhead[2583] = 5'h0d;
assign _c_doomhead[2584] = 5'h08;
assign _c_doomhead[2585] = 5'h02;
assign _c_doomhead[2586] = 5'h08;
assign _c_doomhead[2587] = 5'h00;
assign _c_doomhead[2588] = 5'h00;
assign _c_doomhead[2589] = 5'h00;
assign _c_doomhead[2590] = 5'h00;
assign _c_doomhead[2591] = 5'h00;
assign _c_doomhead[2592] = 5'h00;
assign _c_doomhead[2593] = 5'h00;
assign _c_doomhead[2594] = 5'h00;
assign _c_doomhead[2595] = 5'h01;
assign _c_doomhead[2596] = 5'h02;
assign _c_doomhead[2597] = 5'h01;
assign _c_doomhead[2598] = 5'h0c;
assign _c_doomhead[2599] = 5'h14;
assign _c_doomhead[2600] = 5'h19;
assign _c_doomhead[2601] = 5'h14;
assign _c_doomhead[2602] = 5'h13;
assign _c_doomhead[2603] = 5'h12;
assign _c_doomhead[2604] = 5'h16;
assign _c_doomhead[2605] = 5'h12;
assign _c_doomhead[2606] = 5'h16;
assign _c_doomhead[2607] = 5'h16;
assign _c_doomhead[2608] = 5'h12;
assign _c_doomhead[2609] = 5'h16;
assign _c_doomhead[2610] = 5'h12;
assign _c_doomhead[2611] = 5'h13;
assign _c_doomhead[2612] = 5'h14;
assign _c_doomhead[2613] = 5'h19;
assign _c_doomhead[2614] = 5'h14;
assign _c_doomhead[2615] = 5'h0c;
assign _c_doomhead[2616] = 5'h01;
assign _c_doomhead[2617] = 5'h02;
assign _c_doomhead[2618] = 5'h01;
assign _c_doomhead[2619] = 5'h00;
assign _c_doomhead[2620] = 5'h00;
assign _c_doomhead[2621] = 5'h00;
assign _c_doomhead[2622] = 5'h00;
assign _c_doomhead[2623] = 5'h00;
assign _c_doomhead[2624] = 5'h00;
assign _c_doomhead[2625] = 5'h00;
assign _c_doomhead[2626] = 5'h00;
assign _c_doomhead[2627] = 5'h00;
assign _c_doomhead[2628] = 5'h02;
assign _c_doomhead[2629] = 5'h08;
assign _c_doomhead[2630] = 5'h09;
assign _c_doomhead[2631] = 5'h0b;
assign _c_doomhead[2632] = 5'h0f;
assign _c_doomhead[2633] = 5'h0d;
assign _c_doomhead[2634] = 5'h19;
assign _c_doomhead[2635] = 5'h18;
assign _c_doomhead[2636] = 5'h14;
assign _c_doomhead[2637] = 5'h0d;
assign _c_doomhead[2638] = 5'h18;
assign _c_doomhead[2639] = 5'h16;
assign _c_doomhead[2640] = 5'h0d;
assign _c_doomhead[2641] = 5'h14;
assign _c_doomhead[2642] = 5'h18;
assign _c_doomhead[2643] = 5'h19;
assign _c_doomhead[2644] = 5'h0d;
assign _c_doomhead[2645] = 5'h0f;
assign _c_doomhead[2646] = 5'h0b;
assign _c_doomhead[2647] = 5'h09;
assign _c_doomhead[2648] = 5'h08;
assign _c_doomhead[2649] = 5'h02;
assign _c_doomhead[2650] = 5'h00;
assign _c_doomhead[2651] = 5'h00;
assign _c_doomhead[2652] = 5'h00;
assign _c_doomhead[2653] = 5'h00;
assign _c_doomhead[2654] = 5'h00;
assign _c_doomhead[2655] = 5'h00;
assign _c_doomhead[2656] = 5'h00;
assign _c_doomhead[2657] = 5'h00;
assign _c_doomhead[2658] = 5'h00;
assign _c_doomhead[2659] = 5'h00;
assign _c_doomhead[2660] = 5'h02;
assign _c_doomhead[2661] = 5'h06;
assign _c_doomhead[2662] = 5'h07;
assign _c_doomhead[2663] = 5'h09;
assign _c_doomhead[2664] = 5'h0f;
assign _c_doomhead[2665] = 5'h19;
assign _c_doomhead[2666] = 5'h16;
assign _c_doomhead[2667] = 5'h0d;
assign _c_doomhead[2668] = 5'h0b;
assign _c_doomhead[2669] = 5'h07;
assign _c_doomhead[2670] = 5'h00;
assign _c_doomhead[2671] = 5'h00;
assign _c_doomhead[2672] = 5'h07;
assign _c_doomhead[2673] = 5'h0b;
assign _c_doomhead[2674] = 5'h0d;
assign _c_doomhead[2675] = 5'h16;
assign _c_doomhead[2676] = 5'h19;
assign _c_doomhead[2677] = 5'h0f;
assign _c_doomhead[2678] = 5'h09;
assign _c_doomhead[2679] = 5'h07;
assign _c_doomhead[2680] = 5'h06;
assign _c_doomhead[2681] = 5'h02;
assign _c_doomhead[2682] = 5'h00;
assign _c_doomhead[2683] = 5'h00;
assign _c_doomhead[2684] = 5'h00;
assign _c_doomhead[2685] = 5'h00;
assign _c_doomhead[2686] = 5'h00;
assign _c_doomhead[2687] = 5'h00;
assign _c_doomhead[2688] = 5'h00;
assign _c_doomhead[2689] = 5'h00;
assign _c_doomhead[2690] = 5'h00;
assign _c_doomhead[2691] = 5'h00;
assign _c_doomhead[2692] = 5'h00;
assign _c_doomhead[2693] = 5'h06;
assign _c_doomhead[2694] = 5'h0a;
assign _c_doomhead[2695] = 5'h07;
assign _c_doomhead[2696] = 5'h0d;
assign _c_doomhead[2697] = 5'h16;
assign _c_doomhead[2698] = 5'h12;
assign _c_doomhead[2699] = 5'h09;
assign _c_doomhead[2700] = 5'h0e;
assign _c_doomhead[2701] = 5'h06;
assign _c_doomhead[2702] = 5'h08;
assign _c_doomhead[2703] = 5'h08;
assign _c_doomhead[2704] = 5'h06;
assign _c_doomhead[2705] = 5'h0e;
assign _c_doomhead[2706] = 5'h09;
assign _c_doomhead[2707] = 5'h12;
assign _c_doomhead[2708] = 5'h16;
assign _c_doomhead[2709] = 5'h0d;
assign _c_doomhead[2710] = 5'h07;
assign _c_doomhead[2711] = 5'h0a;
assign _c_doomhead[2712] = 5'h06;
assign _c_doomhead[2713] = 5'h00;
assign _c_doomhead[2714] = 5'h00;
assign _c_doomhead[2715] = 5'h00;
assign _c_doomhead[2716] = 5'h00;
assign _c_doomhead[2717] = 5'h00;
assign _c_doomhead[2718] = 5'h00;
assign _c_doomhead[2719] = 5'h00;
assign _c_doomhead[2720] = 5'h00;
assign _c_doomhead[2721] = 5'h00;
assign _c_doomhead[2722] = 5'h00;
assign _c_doomhead[2723] = 5'h00;
assign _c_doomhead[2724] = 5'h00;
assign _c_doomhead[2725] = 5'h02;
assign _c_doomhead[2726] = 5'h13;
assign _c_doomhead[2727] = 5'h07;
assign _c_doomhead[2728] = 5'h12;
assign _c_doomhead[2729] = 5'h18;
assign _c_doomhead[2730] = 5'h0f;
assign _c_doomhead[2731] = 5'h0c;
assign _c_doomhead[2732] = 5'h14;
assign _c_doomhead[2733] = 5'h0f;
assign _c_doomhead[2734] = 5'h09;
assign _c_doomhead[2735] = 5'h09;
assign _c_doomhead[2736] = 5'h0f;
assign _c_doomhead[2737] = 5'h14;
assign _c_doomhead[2738] = 5'h0c;
assign _c_doomhead[2739] = 5'h0f;
assign _c_doomhead[2740] = 5'h18;
assign _c_doomhead[2741] = 5'h12;
assign _c_doomhead[2742] = 5'h07;
assign _c_doomhead[2743] = 5'h13;
assign _c_doomhead[2744] = 5'h02;
assign _c_doomhead[2745] = 5'h00;
assign _c_doomhead[2746] = 5'h00;
assign _c_doomhead[2747] = 5'h00;
assign _c_doomhead[2748] = 5'h00;
assign _c_doomhead[2749] = 5'h00;
assign _c_doomhead[2750] = 5'h00;
assign _c_doomhead[2751] = 5'h00;
assign _c_doomhead[2752] = 5'h00;
assign _c_doomhead[2753] = 5'h00;
assign _c_doomhead[2754] = 5'h00;
assign _c_doomhead[2755] = 5'h00;
assign _c_doomhead[2756] = 5'h00;
assign _c_doomhead[2757] = 5'h0e;
assign _c_doomhead[2758] = 5'h0b;
assign _c_doomhead[2759] = 5'h09;
assign _c_doomhead[2760] = 5'h0d;
assign _c_doomhead[2761] = 5'h12;
assign _c_doomhead[2762] = 5'h0c;
assign _c_doomhead[2763] = 5'h0d;
assign _c_doomhead[2764] = 5'h18;
assign _c_doomhead[2765] = 5'h16;
assign _c_doomhead[2766] = 5'h0d;
assign _c_doomhead[2767] = 5'h0d;
assign _c_doomhead[2768] = 5'h16;
assign _c_doomhead[2769] = 5'h18;
assign _c_doomhead[2770] = 5'h0d;
assign _c_doomhead[2771] = 5'h0c;
assign _c_doomhead[2772] = 5'h12;
assign _c_doomhead[2773] = 5'h0d;
assign _c_doomhead[2774] = 5'h09;
assign _c_doomhead[2775] = 5'h0b;
assign _c_doomhead[2776] = 5'h0e;
assign _c_doomhead[2777] = 5'h00;
assign _c_doomhead[2778] = 5'h00;
assign _c_doomhead[2779] = 5'h00;
assign _c_doomhead[2780] = 5'h00;
assign _c_doomhead[2781] = 5'h00;
assign _c_doomhead[2782] = 5'h00;
assign _c_doomhead[2783] = 5'h00;
assign _c_doomhead[2784] = 5'h00;
assign _c_doomhead[2785] = 5'h00;
assign _c_doomhead[2786] = 5'h00;
assign _c_doomhead[2787] = 5'h00;
assign _c_doomhead[2788] = 5'h00;
assign _c_doomhead[2789] = 5'h00;
assign _c_doomhead[2790] = 5'h08;
assign _c_doomhead[2791] = 5'h0b;
assign _c_doomhead[2792] = 5'h13;
assign _c_doomhead[2793] = 5'h0d;
assign _c_doomhead[2794] = 5'h01;
assign _c_doomhead[2795] = 5'h06;
assign _c_doomhead[2796] = 5'h1f;
assign _c_doomhead[2797] = 5'h1f;
assign _c_doomhead[2798] = 5'h1f;
assign _c_doomhead[2799] = 5'h1f;
assign _c_doomhead[2800] = 5'h1f;
assign _c_doomhead[2801] = 5'h1f;
assign _c_doomhead[2802] = 5'h06;
assign _c_doomhead[2803] = 5'h01;
assign _c_doomhead[2804] = 5'h0d;
assign _c_doomhead[2805] = 5'h13;
assign _c_doomhead[2806] = 5'h0b;
assign _c_doomhead[2807] = 5'h08;
assign _c_doomhead[2808] = 5'h00;
assign _c_doomhead[2809] = 5'h00;
assign _c_doomhead[2810] = 5'h00;
assign _c_doomhead[2811] = 5'h00;
assign _c_doomhead[2812] = 5'h00;
assign _c_doomhead[2813] = 5'h00;
assign _c_doomhead[2814] = 5'h00;
assign _c_doomhead[2815] = 5'h00;
assign _c_doomhead[2816] = 5'h00;
assign _c_doomhead[2817] = 5'h00;
assign _c_doomhead[2818] = 5'h00;
assign _c_doomhead[2819] = 5'h00;
assign _c_doomhead[2820] = 5'h00;
assign _c_doomhead[2821] = 5'h00;
assign _c_doomhead[2822] = 5'h0e;
assign _c_doomhead[2823] = 5'h01;
assign _c_doomhead[2824] = 5'h0a;
assign _c_doomhead[2825] = 5'h13;
assign _c_doomhead[2826] = 5'h13;
assign _c_doomhead[2827] = 5'h13;
assign _c_doomhead[2828] = 5'h0d;
assign _c_doomhead[2829] = 5'h12;
assign _c_doomhead[2830] = 5'h12;
assign _c_doomhead[2831] = 5'h12;
assign _c_doomhead[2832] = 5'h12;
assign _c_doomhead[2833] = 5'h0d;
assign _c_doomhead[2834] = 5'h13;
assign _c_doomhead[2835] = 5'h13;
assign _c_doomhead[2836] = 5'h13;
assign _c_doomhead[2837] = 5'h0a;
assign _c_doomhead[2838] = 5'h01;
assign _c_doomhead[2839] = 5'h0e;
assign _c_doomhead[2840] = 5'h00;
assign _c_doomhead[2841] = 5'h00;
assign _c_doomhead[2842] = 5'h00;
assign _c_doomhead[2843] = 5'h00;
assign _c_doomhead[2844] = 5'h00;
assign _c_doomhead[2845] = 5'h00;
assign _c_doomhead[2846] = 5'h00;
assign _c_doomhead[2847] = 5'h00;
assign _c_doomhead[2848] = 5'h00;
assign _c_doomhead[2849] = 5'h00;
assign _c_doomhead[2850] = 5'h00;
assign _c_doomhead[2851] = 5'h00;
assign _c_doomhead[2852] = 5'h00;
assign _c_doomhead[2853] = 5'h00;
assign _c_doomhead[2854] = 5'h00;
assign _c_doomhead[2855] = 5'h04;
assign _c_doomhead[2856] = 5'h07;
assign _c_doomhead[2857] = 5'h0c;
assign _c_doomhead[2858] = 5'h14;
assign _c_doomhead[2859] = 5'h13;
assign _c_doomhead[2860] = 5'h0b;
assign _c_doomhead[2861] = 5'h01;
assign _c_doomhead[2862] = 5'h15;
assign _c_doomhead[2863] = 5'h15;
assign _c_doomhead[2864] = 5'h01;
assign _c_doomhead[2865] = 5'h0b;
assign _c_doomhead[2866] = 5'h13;
assign _c_doomhead[2867] = 5'h14;
assign _c_doomhead[2868] = 5'h0c;
assign _c_doomhead[2869] = 5'h07;
assign _c_doomhead[2870] = 5'h04;
assign _c_doomhead[2871] = 5'h00;
assign _c_doomhead[2872] = 5'h00;
assign _c_doomhead[2873] = 5'h00;
assign _c_doomhead[2874] = 5'h00;
assign _c_doomhead[2875] = 5'h00;
assign _c_doomhead[2876] = 5'h00;
assign _c_doomhead[2877] = 5'h00;
assign _c_doomhead[2878] = 5'h00;
assign _c_doomhead[2879] = 5'h00;
assign _c_doomhead[2880] = 5'h00;
assign _c_doomhead[2881] = 5'h00;
assign _c_doomhead[2882] = 5'h00;
assign _c_doomhead[2883] = 5'h00;
assign _c_doomhead[2884] = 5'h00;
assign _c_doomhead[2885] = 5'h00;
assign _c_doomhead[2886] = 5'h00;
assign _c_doomhead[2887] = 5'h00;
assign _c_doomhead[2888] = 5'h04;
assign _c_doomhead[2889] = 5'h09;
assign _c_doomhead[2890] = 5'h0c;
assign _c_doomhead[2891] = 5'h14;
assign _c_doomhead[2892] = 5'h13;
assign _c_doomhead[2893] = 5'h13;
assign _c_doomhead[2894] = 5'h12;
assign _c_doomhead[2895] = 5'h12;
assign _c_doomhead[2896] = 5'h13;
assign _c_doomhead[2897] = 5'h13;
assign _c_doomhead[2898] = 5'h14;
assign _c_doomhead[2899] = 5'h0c;
assign _c_doomhead[2900] = 5'h09;
assign _c_doomhead[2901] = 5'h04;
assign _c_doomhead[2902] = 5'h00;
assign _c_doomhead[2903] = 5'h00;
assign _c_doomhead[2904] = 5'h00;
assign _c_doomhead[2905] = 5'h00;
assign _c_doomhead[2906] = 5'h00;
assign _c_doomhead[2907] = 5'h00;
assign _c_doomhead[2908] = 5'h00;
assign _c_doomhead[2909] = 5'h00;
assign _c_doomhead[2910] = 5'h00;
assign _c_doomhead[2911] = 5'h00;
assign _c_doomhead[2912] = 5'h00;
assign _c_doomhead[2913] = 5'h00;
assign _c_doomhead[2914] = 5'h00;
assign _c_doomhead[2915] = 5'h00;
assign _c_doomhead[2916] = 5'h00;
assign _c_doomhead[2917] = 5'h00;
assign _c_doomhead[2918] = 5'h00;
assign _c_doomhead[2919] = 5'h00;
assign _c_doomhead[2920] = 5'h00;
assign _c_doomhead[2921] = 5'h0e;
assign _c_doomhead[2922] = 5'h08;
assign _c_doomhead[2923] = 5'h0a;
assign _c_doomhead[2924] = 5'h0d;
assign _c_doomhead[2925] = 5'h12;
assign _c_doomhead[2926] = 5'h16;
assign _c_doomhead[2927] = 5'h16;
assign _c_doomhead[2928] = 5'h12;
assign _c_doomhead[2929] = 5'h0d;
assign _c_doomhead[2930] = 5'h0a;
assign _c_doomhead[2931] = 5'h08;
assign _c_doomhead[2932] = 5'h0e;
assign _c_doomhead[2933] = 5'h00;
assign _c_doomhead[2934] = 5'h00;
assign _c_doomhead[2935] = 5'h00;
assign _c_doomhead[2936] = 5'h00;
assign _c_doomhead[2937] = 5'h00;
assign _c_doomhead[2938] = 5'h00;
assign _c_doomhead[2939] = 5'h00;
assign _c_doomhead[2940] = 5'h00;
assign _c_doomhead[2941] = 5'h00;
assign _c_doomhead[2942] = 5'h00;
assign _c_doomhead[2943] = 5'h00;
assign _c_doomhead[2944] = 5'h00;
assign _c_doomhead[2945] = 5'h00;
assign _c_doomhead[2946] = 5'h00;
assign _c_doomhead[2947] = 5'h00;
assign _c_doomhead[2948] = 5'h00;
assign _c_doomhead[2949] = 5'h00;
assign _c_doomhead[2950] = 5'h00;
assign _c_doomhead[2951] = 5'h00;
assign _c_doomhead[2952] = 5'h00;
assign _c_doomhead[2953] = 5'h00;
assign _c_doomhead[2954] = 5'h00;
assign _c_doomhead[2955] = 5'h04;
assign _c_doomhead[2956] = 5'h01;
assign _c_doomhead[2957] = 5'h09;
assign _c_doomhead[2958] = 5'h09;
assign _c_doomhead[2959] = 5'h09;
assign _c_doomhead[2960] = 5'h09;
assign _c_doomhead[2961] = 5'h01;
assign _c_doomhead[2962] = 5'h04;
assign _c_doomhead[2963] = 5'h00;
assign _c_doomhead[2964] = 5'h00;
assign _c_doomhead[2965] = 5'h00;
assign _c_doomhead[2966] = 5'h00;
assign _c_doomhead[2967] = 5'h00;
assign _c_doomhead[2968] = 5'h00;
assign _c_doomhead[2969] = 5'h00;
assign _c_doomhead[2970] = 5'h00;
assign _c_doomhead[2971] = 5'h00;
assign _c_doomhead[2972] = 5'h00;
assign _c_doomhead[2973] = 5'h00;
assign _c_doomhead[2974] = 5'h00;
assign _c_doomhead[2975] = 5'h00;
assign _c_doomhead[2976] = 5'h00;
assign _c_doomhead[2977] = 5'h00;
assign _c_doomhead[2978] = 5'h00;
assign _c_doomhead[2979] = 5'h00;
assign _c_doomhead[2980] = 5'h00;
assign _c_doomhead[2981] = 5'h00;
assign _c_doomhead[2982] = 5'h00;
assign _c_doomhead[2983] = 5'h00;
assign _c_doomhead[2984] = 5'h00;
assign _c_doomhead[2985] = 5'h00;
assign _c_doomhead[2986] = 5'h00;
assign _c_doomhead[2987] = 5'h00;
assign _c_doomhead[2988] = 5'h00;
assign _c_doomhead[2989] = 5'h00;
assign _c_doomhead[2990] = 5'h00;
assign _c_doomhead[2991] = 5'h00;
assign _c_doomhead[2992] = 5'h00;
assign _c_doomhead[2993] = 5'h00;
assign _c_doomhead[2994] = 5'h00;
assign _c_doomhead[2995] = 5'h00;
assign _c_doomhead[2996] = 5'h00;
assign _c_doomhead[2997] = 5'h00;
assign _c_doomhead[2998] = 5'h00;
assign _c_doomhead[2999] = 5'h00;
assign _c_doomhead[3000] = 5'h00;
assign _c_doomhead[3001] = 5'h00;
assign _c_doomhead[3002] = 5'h00;
assign _c_doomhead[3003] = 5'h00;
assign _c_doomhead[3004] = 5'h00;
assign _c_doomhead[3005] = 5'h00;
assign _c_doomhead[3006] = 5'h00;
assign _c_doomhead[3007] = 5'h00;
assign _c_doomhead[3008] = 5'h00;
assign _c_doomhead[3009] = 5'h00;
assign _c_doomhead[3010] = 5'h00;
assign _c_doomhead[3011] = 5'h00;
assign _c_doomhead[3012] = 5'h00;
assign _c_doomhead[3013] = 5'h00;
assign _c_doomhead[3014] = 5'h00;
assign _c_doomhead[3015] = 5'h00;
assign _c_doomhead[3016] = 5'h00;
assign _c_doomhead[3017] = 5'h00;
assign _c_doomhead[3018] = 5'h00;
assign _c_doomhead[3019] = 5'h00;
assign _c_doomhead[3020] = 5'h00;
assign _c_doomhead[3021] = 5'h00;
assign _c_doomhead[3022] = 5'h00;
assign _c_doomhead[3023] = 5'h00;
assign _c_doomhead[3024] = 5'h00;
assign _c_doomhead[3025] = 5'h00;
assign _c_doomhead[3026] = 5'h00;
assign _c_doomhead[3027] = 5'h00;
assign _c_doomhead[3028] = 5'h00;
assign _c_doomhead[3029] = 5'h00;
assign _c_doomhead[3030] = 5'h00;
assign _c_doomhead[3031] = 5'h00;
assign _c_doomhead[3032] = 5'h00;
assign _c_doomhead[3033] = 5'h00;
assign _c_doomhead[3034] = 5'h00;
assign _c_doomhead[3035] = 5'h00;
assign _c_doomhead[3036] = 5'h00;
assign _c_doomhead[3037] = 5'h00;
assign _c_doomhead[3038] = 5'h00;
assign _c_doomhead[3039] = 5'h00;
assign _c_doomhead[3040] = 5'h00;
assign _c_doomhead[3041] = 5'h00;
assign _c_doomhead[3042] = 5'h00;
assign _c_doomhead[3043] = 5'h00;
assign _c_doomhead[3044] = 5'h00;
assign _c_doomhead[3045] = 5'h00;
assign _c_doomhead[3046] = 5'h00;
assign _c_doomhead[3047] = 5'h00;
assign _c_doomhead[3048] = 5'h00;
assign _c_doomhead[3049] = 5'h00;
assign _c_doomhead[3050] = 5'h00;
assign _c_doomhead[3051] = 5'h00;
assign _c_doomhead[3052] = 5'h00;
assign _c_doomhead[3053] = 5'h00;
assign _c_doomhead[3054] = 5'h00;
assign _c_doomhead[3055] = 5'h00;
assign _c_doomhead[3056] = 5'h00;
assign _c_doomhead[3057] = 5'h00;
assign _c_doomhead[3058] = 5'h00;
assign _c_doomhead[3059] = 5'h00;
assign _c_doomhead[3060] = 5'h00;
assign _c_doomhead[3061] = 5'h00;
assign _c_doomhead[3062] = 5'h00;
assign _c_doomhead[3063] = 5'h00;
assign _c_doomhead[3064] = 5'h00;
assign _c_doomhead[3065] = 5'h00;
assign _c_doomhead[3066] = 5'h00;
assign _c_doomhead[3067] = 5'h00;
assign _c_doomhead[3068] = 5'h00;
assign _c_doomhead[3069] = 5'h00;
assign _c_doomhead[3070] = 5'h00;
assign _c_doomhead[3071] = 5'h00;
assign _c_doomhead[3072] = 5'h00;
assign _c_doomhead[3073] = 5'h00;
assign _c_doomhead[3074] = 5'h00;
assign _c_doomhead[3075] = 5'h00;
assign _c_doomhead[3076] = 5'h00;
assign _c_doomhead[3077] = 5'h00;
assign _c_doomhead[3078] = 5'h00;
assign _c_doomhead[3079] = 5'h00;
assign _c_doomhead[3080] = 5'h00;
assign _c_doomhead[3081] = 5'h00;
assign _c_doomhead[3082] = 5'h00;
assign _c_doomhead[3083] = 5'h03;
assign _c_doomhead[3084] = 5'h03;
assign _c_doomhead[3085] = 5'h03;
assign _c_doomhead[3086] = 5'h03;
assign _c_doomhead[3087] = 5'h03;
assign _c_doomhead[3088] = 5'h03;
assign _c_doomhead[3089] = 5'h03;
assign _c_doomhead[3090] = 5'h03;
assign _c_doomhead[3091] = 5'h05;
assign _c_doomhead[3092] = 5'h05;
assign _c_doomhead[3093] = 5'h05;
assign _c_doomhead[3094] = 5'h00;
assign _c_doomhead[3095] = 5'h00;
assign _c_doomhead[3096] = 5'h00;
assign _c_doomhead[3097] = 5'h00;
assign _c_doomhead[3098] = 5'h00;
assign _c_doomhead[3099] = 5'h00;
assign _c_doomhead[3100] = 5'h00;
assign _c_doomhead[3101] = 5'h00;
assign _c_doomhead[3102] = 5'h00;
assign _c_doomhead[3103] = 5'h00;
assign _c_doomhead[3104] = 5'h00;
assign _c_doomhead[3105] = 5'h00;
assign _c_doomhead[3106] = 5'h00;
assign _c_doomhead[3107] = 5'h00;
assign _c_doomhead[3108] = 5'h00;
assign _c_doomhead[3109] = 5'h00;
assign _c_doomhead[3110] = 5'h00;
assign _c_doomhead[3111] = 5'h00;
assign _c_doomhead[3112] = 5'h03;
assign _c_doomhead[3113] = 5'h03;
assign _c_doomhead[3114] = 5'h02;
assign _c_doomhead[3115] = 5'h02;
assign _c_doomhead[3116] = 5'h04;
assign _c_doomhead[3117] = 5'h08;
assign _c_doomhead[3118] = 5'h08;
assign _c_doomhead[3119] = 5'h08;
assign _c_doomhead[3120] = 5'h06;
assign _c_doomhead[3121] = 5'h06;
assign _c_doomhead[3122] = 5'h04;
assign _c_doomhead[3123] = 5'h04;
assign _c_doomhead[3124] = 5'h02;
assign _c_doomhead[3125] = 5'h05;
assign _c_doomhead[3126] = 5'h05;
assign _c_doomhead[3127] = 5'h05;
assign _c_doomhead[3128] = 5'h00;
assign _c_doomhead[3129] = 5'h00;
assign _c_doomhead[3130] = 5'h00;
assign _c_doomhead[3131] = 5'h00;
assign _c_doomhead[3132] = 5'h00;
assign _c_doomhead[3133] = 5'h00;
assign _c_doomhead[3134] = 5'h00;
assign _c_doomhead[3135] = 5'h00;
assign _c_doomhead[3136] = 5'h00;
assign _c_doomhead[3137] = 5'h00;
assign _c_doomhead[3138] = 5'h00;
assign _c_doomhead[3139] = 5'h00;
assign _c_doomhead[3140] = 5'h00;
assign _c_doomhead[3141] = 5'h00;
assign _c_doomhead[3142] = 5'h00;
assign _c_doomhead[3143] = 5'h05;
assign _c_doomhead[3144] = 5'h02;
assign _c_doomhead[3145] = 5'h04;
assign _c_doomhead[3146] = 5'h08;
assign _c_doomhead[3147] = 5'h01;
assign _c_doomhead[3148] = 5'h0a;
assign _c_doomhead[3149] = 5'h0a;
assign _c_doomhead[3150] = 5'h07;
assign _c_doomhead[3151] = 5'h07;
assign _c_doomhead[3152] = 5'h01;
assign _c_doomhead[3153] = 5'h08;
assign _c_doomhead[3154] = 5'h06;
assign _c_doomhead[3155] = 5'h04;
assign _c_doomhead[3156] = 5'h02;
assign _c_doomhead[3157] = 5'h05;
assign _c_doomhead[3158] = 5'h05;
assign _c_doomhead[3159] = 5'h05;
assign _c_doomhead[3160] = 5'h03;
assign _c_doomhead[3161] = 5'h03;
assign _c_doomhead[3162] = 5'h00;
assign _c_doomhead[3163] = 5'h00;
assign _c_doomhead[3164] = 5'h00;
assign _c_doomhead[3165] = 5'h00;
assign _c_doomhead[3166] = 5'h00;
assign _c_doomhead[3167] = 5'h00;
assign _c_doomhead[3168] = 5'h00;
assign _c_doomhead[3169] = 5'h00;
assign _c_doomhead[3170] = 5'h00;
assign _c_doomhead[3171] = 5'h00;
assign _c_doomhead[3172] = 5'h00;
assign _c_doomhead[3173] = 5'h05;
assign _c_doomhead[3174] = 5'h03;
assign _c_doomhead[3175] = 5'h05;
assign _c_doomhead[3176] = 5'h02;
assign _c_doomhead[3177] = 5'h04;
assign _c_doomhead[3178] = 5'h08;
assign _c_doomhead[3179] = 5'h01;
assign _c_doomhead[3180] = 5'h07;
assign _c_doomhead[3181] = 5'h07;
assign _c_doomhead[3182] = 5'h07;
assign _c_doomhead[3183] = 5'h07;
assign _c_doomhead[3184] = 5'h01;
assign _c_doomhead[3185] = 5'h08;
assign _c_doomhead[3186] = 5'h06;
assign _c_doomhead[3187] = 5'h02;
assign _c_doomhead[3188] = 5'h02;
assign _c_doomhead[3189] = 5'h05;
assign _c_doomhead[3190] = 5'h05;
assign _c_doomhead[3191] = 5'h10;
assign _c_doomhead[3192] = 5'h10;
assign _c_doomhead[3193] = 5'h03;
assign _c_doomhead[3194] = 5'h03;
assign _c_doomhead[3195] = 5'h00;
assign _c_doomhead[3196] = 5'h00;
assign _c_doomhead[3197] = 5'h00;
assign _c_doomhead[3198] = 5'h00;
assign _c_doomhead[3199] = 5'h00;
assign _c_doomhead[3200] = 5'h00;
assign _c_doomhead[3201] = 5'h00;
assign _c_doomhead[3202] = 5'h00;
assign _c_doomhead[3203] = 5'h00;
assign _c_doomhead[3204] = 5'h05;
assign _c_doomhead[3205] = 5'h05;
assign _c_doomhead[3206] = 5'h05;
assign _c_doomhead[3207] = 5'h02;
assign _c_doomhead[3208] = 5'h01;
assign _c_doomhead[3209] = 5'h0a;
assign _c_doomhead[3210] = 5'h0f;
assign _c_doomhead[3211] = 5'h0f;
assign _c_doomhead[3212] = 5'h0a;
assign _c_doomhead[3213] = 5'h07;
assign _c_doomhead[3214] = 5'h01;
assign _c_doomhead[3215] = 5'h08;
assign _c_doomhead[3216] = 5'h06;
assign _c_doomhead[3217] = 5'h02;
assign _c_doomhead[3218] = 5'h02;
assign _c_doomhead[3219] = 5'h02;
assign _c_doomhead[3220] = 5'h05;
assign _c_doomhead[3221] = 5'h05;
assign _c_doomhead[3222] = 5'h10;
assign _c_doomhead[3223] = 5'h05;
assign _c_doomhead[3224] = 5'h03;
assign _c_doomhead[3225] = 5'h10;
assign _c_doomhead[3226] = 5'h03;
assign _c_doomhead[3227] = 5'h03;
assign _c_doomhead[3228] = 5'h00;
assign _c_doomhead[3229] = 5'h00;
assign _c_doomhead[3230] = 5'h00;
assign _c_doomhead[3231] = 5'h00;
assign _c_doomhead[3232] = 5'h00;
assign _c_doomhead[3233] = 5'h00;
assign _c_doomhead[3234] = 5'h00;
assign _c_doomhead[3235] = 5'h02;
assign _c_doomhead[3236] = 5'h05;
assign _c_doomhead[3237] = 5'h05;
assign _c_doomhead[3238] = 5'h02;
assign _c_doomhead[3239] = 5'h01;
assign _c_doomhead[3240] = 5'h07;
assign _c_doomhead[3241] = 5'h07;
assign _c_doomhead[3242] = 5'h07;
assign _c_doomhead[3243] = 5'h07;
assign _c_doomhead[3244] = 5'h07;
assign _c_doomhead[3245] = 5'h01;
assign _c_doomhead[3246] = 5'h08;
assign _c_doomhead[3247] = 5'h06;
assign _c_doomhead[3248] = 5'h02;
assign _c_doomhead[3249] = 5'h02;
assign _c_doomhead[3250] = 5'h02;
assign _c_doomhead[3251] = 5'h02;
assign _c_doomhead[3252] = 5'h05;
assign _c_doomhead[3253] = 5'h05;
assign _c_doomhead[3254] = 5'h10;
assign _c_doomhead[3255] = 5'h10;
assign _c_doomhead[3256] = 5'h05;
assign _c_doomhead[3257] = 5'h10;
assign _c_doomhead[3258] = 5'h03;
assign _c_doomhead[3259] = 5'h03;
assign _c_doomhead[3260] = 5'h00;
assign _c_doomhead[3261] = 5'h00;
assign _c_doomhead[3262] = 5'h00;
assign _c_doomhead[3263] = 5'h00;
assign _c_doomhead[3264] = 5'h00;
assign _c_doomhead[3265] = 5'h00;
assign _c_doomhead[3266] = 5'h05;
assign _c_doomhead[3267] = 5'h02;
assign _c_doomhead[3268] = 5'h06;
assign _c_doomhead[3269] = 5'h06;
assign _c_doomhead[3270] = 5'h04;
assign _c_doomhead[3271] = 5'h06;
assign _c_doomhead[3272] = 5'h06;
assign _c_doomhead[3273] = 5'h06;
assign _c_doomhead[3274] = 5'h06;
assign _c_doomhead[3275] = 5'h01;
assign _c_doomhead[3276] = 5'h01;
assign _c_doomhead[3277] = 5'h06;
assign _c_doomhead[3278] = 5'h06;
assign _c_doomhead[3279] = 5'h04;
assign _c_doomhead[3280] = 5'h02;
assign _c_doomhead[3281] = 5'h02;
assign _c_doomhead[3282] = 5'h02;
assign _c_doomhead[3283] = 5'h05;
assign _c_doomhead[3284] = 5'h05;
assign _c_doomhead[3285] = 5'h05;
assign _c_doomhead[3286] = 5'h05;
assign _c_doomhead[3287] = 5'h10;
assign _c_doomhead[3288] = 5'h10;
assign _c_doomhead[3289] = 5'h10;
assign _c_doomhead[3290] = 5'h10;
assign _c_doomhead[3291] = 5'h03;
assign _c_doomhead[3292] = 5'h03;
assign _c_doomhead[3293] = 5'h00;
assign _c_doomhead[3294] = 5'h00;
assign _c_doomhead[3295] = 5'h00;
assign _c_doomhead[3296] = 5'h00;
assign _c_doomhead[3297] = 5'h11;
assign _c_doomhead[3298] = 5'h04;
assign _c_doomhead[3299] = 5'h08;
assign _c_doomhead[3300] = 5'h07;
assign _c_doomhead[3301] = 5'h08;
assign _c_doomhead[3302] = 5'h08;
assign _c_doomhead[3303] = 5'h01;
assign _c_doomhead[3304] = 5'h01;
assign _c_doomhead[3305] = 5'h06;
assign _c_doomhead[3306] = 5'h04;
assign _c_doomhead[3307] = 5'h04;
assign _c_doomhead[3308] = 5'h04;
assign _c_doomhead[3309] = 5'h01;
assign _c_doomhead[3310] = 5'h09;
assign _c_doomhead[3311] = 5'h02;
assign _c_doomhead[3312] = 5'h0e;
assign _c_doomhead[3313] = 5'h0e;
assign _c_doomhead[3314] = 5'h04;
assign _c_doomhead[3315] = 5'h0e;
assign _c_doomhead[3316] = 5'h10;
assign _c_doomhead[3317] = 5'h10;
assign _c_doomhead[3318] = 5'h05;
assign _c_doomhead[3319] = 5'h05;
assign _c_doomhead[3320] = 5'h10;
assign _c_doomhead[3321] = 5'h10;
assign _c_doomhead[3322] = 5'h10;
assign _c_doomhead[3323] = 5'h03;
assign _c_doomhead[3324] = 5'h03;
assign _c_doomhead[3325] = 5'h00;
assign _c_doomhead[3326] = 5'h00;
assign _c_doomhead[3327] = 5'h00;
assign _c_doomhead[3328] = 5'h00;
assign _c_doomhead[3329] = 5'h11;
assign _c_doomhead[3330] = 5'h10;
assign _c_doomhead[3331] = 5'h10;
assign _c_doomhead[3332] = 5'h10;
assign _c_doomhead[3333] = 5'h07;
assign _c_doomhead[3334] = 5'h08;
assign _c_doomhead[3335] = 5'h04;
assign _c_doomhead[3336] = 5'h02;
assign _c_doomhead[3337] = 5'h04;
assign _c_doomhead[3338] = 5'h06;
assign _c_doomhead[3339] = 5'h05;
assign _c_doomhead[3340] = 5'h05;
assign _c_doomhead[3341] = 5'h02;
assign _c_doomhead[3342] = 5'h02;
assign _c_doomhead[3343] = 5'h15;
assign _c_doomhead[3344] = 5'h01;
assign _c_doomhead[3345] = 5'h04;
assign _c_doomhead[3346] = 5'h0e;
assign _c_doomhead[3347] = 5'h04;
assign _c_doomhead[3348] = 5'h04;
assign _c_doomhead[3349] = 5'h05;
assign _c_doomhead[3350] = 5'h10;
assign _c_doomhead[3351] = 5'h03;
assign _c_doomhead[3352] = 5'h05;
assign _c_doomhead[3353] = 5'h03;
assign _c_doomhead[3354] = 5'h03;
assign _c_doomhead[3355] = 5'h10;
assign _c_doomhead[3356] = 5'h03;
assign _c_doomhead[3357] = 5'h03;
assign _c_doomhead[3358] = 5'h00;
assign _c_doomhead[3359] = 5'h00;
assign _c_doomhead[3360] = 5'h11;
assign _c_doomhead[3361] = 5'h05;
assign _c_doomhead[3362] = 5'h11;
assign _c_doomhead[3363] = 5'h11;
assign _c_doomhead[3364] = 5'h11;
assign _c_doomhead[3365] = 5'h02;
assign _c_doomhead[3366] = 5'h04;
assign _c_doomhead[3367] = 5'h07;
assign _c_doomhead[3368] = 5'h04;
assign _c_doomhead[3369] = 5'h04;
assign _c_doomhead[3370] = 5'h05;
assign _c_doomhead[3371] = 5'h04;
assign _c_doomhead[3372] = 5'h05;
assign _c_doomhead[3373] = 5'h10;
assign _c_doomhead[3374] = 5'h03;
assign _c_doomhead[3375] = 5'h10;
assign _c_doomhead[3376] = 5'h10;
assign _c_doomhead[3377] = 5'h04;
assign _c_doomhead[3378] = 5'h01;
assign _c_doomhead[3379] = 5'h02;
assign _c_doomhead[3380] = 5'h05;
assign _c_doomhead[3381] = 5'h04;
assign _c_doomhead[3382] = 5'h05;
assign _c_doomhead[3383] = 5'h10;
assign _c_doomhead[3384] = 5'h03;
assign _c_doomhead[3385] = 5'h03;
assign _c_doomhead[3386] = 5'h03;
assign _c_doomhead[3387] = 5'h10;
assign _c_doomhead[3388] = 5'h03;
assign _c_doomhead[3389] = 5'h03;
assign _c_doomhead[3390] = 5'h00;
assign _c_doomhead[3391] = 5'h00;
assign _c_doomhead[3392] = 5'h11;
assign _c_doomhead[3393] = 5'h11;
assign _c_doomhead[3394] = 5'h11;
assign _c_doomhead[3395] = 5'h11;
assign _c_doomhead[3396] = 5'h11;
assign _c_doomhead[3397] = 5'h11;
assign _c_doomhead[3398] = 5'h02;
assign _c_doomhead[3399] = 5'h05;
assign _c_doomhead[3400] = 5'h05;
assign _c_doomhead[3401] = 5'h11;
assign _c_doomhead[3402] = 5'h11;
assign _c_doomhead[3403] = 5'h03;
assign _c_doomhead[3404] = 5'h04;
assign _c_doomhead[3405] = 5'h0e;
assign _c_doomhead[3406] = 5'h06;
assign _c_doomhead[3407] = 5'h06;
assign _c_doomhead[3408] = 5'h02;
assign _c_doomhead[3409] = 5'h03;
assign _c_doomhead[3410] = 5'h02;
assign _c_doomhead[3411] = 5'h06;
assign _c_doomhead[3412] = 5'h02;
assign _c_doomhead[3413] = 5'h05;
assign _c_doomhead[3414] = 5'h04;
assign _c_doomhead[3415] = 5'h05;
assign _c_doomhead[3416] = 5'h10;
assign _c_doomhead[3417] = 5'h03;
assign _c_doomhead[3418] = 5'h03;
assign _c_doomhead[3419] = 5'h10;
assign _c_doomhead[3420] = 5'h03;
assign _c_doomhead[3421] = 5'h03;
assign _c_doomhead[3422] = 5'h00;
assign _c_doomhead[3423] = 5'h00;
assign _c_doomhead[3424] = 5'h00;
assign _c_doomhead[3425] = 5'h11;
assign _c_doomhead[3426] = 5'h05;
assign _c_doomhead[3427] = 5'h02;
assign _c_doomhead[3428] = 5'h11;
assign _c_doomhead[3429] = 5'h1c;
assign _c_doomhead[3430] = 5'h01;
assign _c_doomhead[3431] = 5'h01;
assign _c_doomhead[3432] = 5'h0e;
assign _c_doomhead[3433] = 5'h11;
assign _c_doomhead[3434] = 5'h1b;
assign _c_doomhead[3435] = 5'h1a;
assign _c_doomhead[3436] = 5'h03;
assign _c_doomhead[3437] = 5'h04;
assign _c_doomhead[3438] = 5'h01;
assign _c_doomhead[3439] = 5'h09;
assign _c_doomhead[3440] = 5'h07;
assign _c_doomhead[3441] = 5'h02;
assign _c_doomhead[3442] = 5'h03;
assign _c_doomhead[3443] = 5'h02;
assign _c_doomhead[3444] = 5'h06;
assign _c_doomhead[3445] = 5'h02;
assign _c_doomhead[3446] = 5'h05;
assign _c_doomhead[3447] = 5'h0e;
assign _c_doomhead[3448] = 5'h10;
assign _c_doomhead[3449] = 5'h03;
assign _c_doomhead[3450] = 5'h03;
assign _c_doomhead[3451] = 5'h10;
assign _c_doomhead[3452] = 5'h03;
assign _c_doomhead[3453] = 5'h03;
assign _c_doomhead[3454] = 5'h00;
assign _c_doomhead[3455] = 5'h00;
assign _c_doomhead[3456] = 5'h00;
assign _c_doomhead[3457] = 5'h00;
assign _c_doomhead[3458] = 5'h05;
assign _c_doomhead[3459] = 5'h01;
assign _c_doomhead[3460] = 5'h1c;
assign _c_doomhead[3461] = 5'h1c;
assign _c_doomhead[3462] = 5'h0d;
assign _c_doomhead[3463] = 5'h0d;
assign _c_doomhead[3464] = 5'h09;
assign _c_doomhead[3465] = 5'h0e;
assign _c_doomhead[3466] = 5'h1a;
assign _c_doomhead[3467] = 5'h1a;
assign _c_doomhead[3468] = 5'h1a;
assign _c_doomhead[3469] = 5'h04;
assign _c_doomhead[3470] = 5'h08;
assign _c_doomhead[3471] = 5'h0b;
assign _c_doomhead[3472] = 5'h01;
assign _c_doomhead[3473] = 5'h07;
assign _c_doomhead[3474] = 5'h0e;
assign _c_doomhead[3475] = 5'h05;
assign _c_doomhead[3476] = 5'h02;
assign _c_doomhead[3477] = 5'h05;
assign _c_doomhead[3478] = 5'h03;
assign _c_doomhead[3479] = 5'h03;
assign _c_doomhead[3480] = 5'h0e;
assign _c_doomhead[3481] = 5'h10;
assign _c_doomhead[3482] = 5'h03;
assign _c_doomhead[3483] = 5'h03;
assign _c_doomhead[3484] = 5'h03;
assign _c_doomhead[3485] = 5'h03;
assign _c_doomhead[3486] = 5'h00;
assign _c_doomhead[3487] = 5'h00;
assign _c_doomhead[3488] = 5'h00;
assign _c_doomhead[3489] = 5'h00;
assign _c_doomhead[3490] = 5'h00;
assign _c_doomhead[3491] = 5'h09;
assign _c_doomhead[3492] = 5'h1c;
assign _c_doomhead[3493] = 5'h1c;
assign _c_doomhead[3494] = 5'h0d;
assign _c_doomhead[3495] = 5'h0d;
assign _c_doomhead[3496] = 5'h0d;
assign _c_doomhead[3497] = 5'h0d;
assign _c_doomhead[3498] = 5'h0e;
assign _c_doomhead[3499] = 5'h1a;
assign _c_doomhead[3500] = 5'h1d;
assign _c_doomhead[3501] = 5'h0d;
assign _c_doomhead[3502] = 5'h0b;
assign _c_doomhead[3503] = 5'h0b;
assign _c_doomhead[3504] = 5'h01;
assign _c_doomhead[3505] = 5'h01;
assign _c_doomhead[3506] = 5'h15;
assign _c_doomhead[3507] = 5'h05;
assign _c_doomhead[3508] = 5'h05;
assign _c_doomhead[3509] = 5'h04;
assign _c_doomhead[3510] = 5'h04;
assign _c_doomhead[3511] = 5'h04;
assign _c_doomhead[3512] = 5'h04;
assign _c_doomhead[3513] = 5'h0e;
assign _c_doomhead[3514] = 5'h03;
assign _c_doomhead[3515] = 5'h03;
assign _c_doomhead[3516] = 5'h03;
assign _c_doomhead[3517] = 5'h03;
assign _c_doomhead[3518] = 5'h00;
assign _c_doomhead[3519] = 5'h00;
assign _c_doomhead[3520] = 5'h00;
assign _c_doomhead[3521] = 5'h00;
assign _c_doomhead[3522] = 5'h00;
assign _c_doomhead[3523] = 5'h0b;
assign _c_doomhead[3524] = 5'h1a;
assign _c_doomhead[3525] = 5'h1c;
assign _c_doomhead[3526] = 5'h1e;
assign _c_doomhead[3527] = 5'h0d;
assign _c_doomhead[3528] = 5'h19;
assign _c_doomhead[3529] = 5'h18;
assign _c_doomhead[3530] = 5'h18;
assign _c_doomhead[3531] = 5'h1d;
assign _c_doomhead[3532] = 5'h1e;
assign _c_doomhead[3533] = 5'h19;
assign _c_doomhead[3534] = 5'h14;
assign _c_doomhead[3535] = 5'h0f;
assign _c_doomhead[3536] = 5'h0b;
assign _c_doomhead[3537] = 5'h01;
assign _c_doomhead[3538] = 5'h15;
assign _c_doomhead[3539] = 5'h04;
assign _c_doomhead[3540] = 5'h04;
assign _c_doomhead[3541] = 5'h01;
assign _c_doomhead[3542] = 5'h02;
assign _c_doomhead[3543] = 5'h07;
assign _c_doomhead[3544] = 5'h08;
assign _c_doomhead[3545] = 5'h08;
assign _c_doomhead[3546] = 5'h03;
assign _c_doomhead[3547] = 5'h03;
assign _c_doomhead[3548] = 5'h03;
assign _c_doomhead[3549] = 5'h03;
assign _c_doomhead[3550] = 5'h00;
assign _c_doomhead[3551] = 5'h00;
assign _c_doomhead[3552] = 5'h00;
assign _c_doomhead[3553] = 5'h00;
assign _c_doomhead[3554] = 5'h00;
assign _c_doomhead[3555] = 5'h02;
assign _c_doomhead[3556] = 5'h1b;
assign _c_doomhead[3557] = 5'h1a;
assign _c_doomhead[3558] = 5'h1e;
assign _c_doomhead[3559] = 5'h16;
assign _c_doomhead[3560] = 5'h16;
assign _c_doomhead[3561] = 5'h16;
assign _c_doomhead[3562] = 5'h16;
assign _c_doomhead[3563] = 5'h1e;
assign _c_doomhead[3564] = 5'h1e;
assign _c_doomhead[3565] = 5'h16;
assign _c_doomhead[3566] = 5'h18;
assign _c_doomhead[3567] = 5'h14;
assign _c_doomhead[3568] = 5'h0c;
assign _c_doomhead[3569] = 5'h0b;
assign _c_doomhead[3570] = 5'h01;
assign _c_doomhead[3571] = 5'h01;
assign _c_doomhead[3572] = 5'h01;
assign _c_doomhead[3573] = 5'h07;
assign _c_doomhead[3574] = 5'h07;
assign _c_doomhead[3575] = 5'h08;
assign _c_doomhead[3576] = 5'h0a;
assign _c_doomhead[3577] = 5'h08;
assign _c_doomhead[3578] = 5'h03;
assign _c_doomhead[3579] = 5'h03;
assign _c_doomhead[3580] = 5'h03;
assign _c_doomhead[3581] = 5'h03;
assign _c_doomhead[3582] = 5'h00;
assign _c_doomhead[3583] = 5'h00;
assign _c_doomhead[3584] = 5'h00;
assign _c_doomhead[3585] = 5'h00;
assign _c_doomhead[3586] = 5'h00;
assign _c_doomhead[3587] = 5'h10;
assign _c_doomhead[3588] = 5'h10;
assign _c_doomhead[3589] = 5'h02;
assign _c_doomhead[3590] = 5'h0b;
assign _c_doomhead[3591] = 5'h0c;
assign _c_doomhead[3592] = 5'h14;
assign _c_doomhead[3593] = 5'h0f;
assign _c_doomhead[3594] = 5'h07;
assign _c_doomhead[3595] = 5'h04;
assign _c_doomhead[3596] = 5'h04;
assign _c_doomhead[3597] = 5'h09;
assign _c_doomhead[3598] = 5'h0f;
assign _c_doomhead[3599] = 5'h12;
assign _c_doomhead[3600] = 5'h0d;
assign _c_doomhead[3601] = 5'h0c;
assign _c_doomhead[3602] = 5'h09;
assign _c_doomhead[3603] = 5'h09;
assign _c_doomhead[3604] = 5'h09;
assign _c_doomhead[3605] = 5'h09;
assign _c_doomhead[3606] = 5'h0f;
assign _c_doomhead[3607] = 5'h0e;
assign _c_doomhead[3608] = 5'h0a;
assign _c_doomhead[3609] = 5'h01;
assign _c_doomhead[3610] = 5'h03;
assign _c_doomhead[3611] = 5'h03;
assign _c_doomhead[3612] = 5'h03;
assign _c_doomhead[3613] = 5'h03;
assign _c_doomhead[3614] = 5'h00;
assign _c_doomhead[3615] = 5'h00;
assign _c_doomhead[3616] = 5'h00;
assign _c_doomhead[3617] = 5'h00;
assign _c_doomhead[3618] = 5'h00;
assign _c_doomhead[3619] = 5'h00;
assign _c_doomhead[3620] = 5'h10;
assign _c_doomhead[3621] = 5'h17;
assign _c_doomhead[3622] = 5'h1a;
assign _c_doomhead[3623] = 5'h17;
assign _c_doomhead[3624] = 5'h0b;
assign _c_doomhead[3625] = 5'h05;
assign _c_doomhead[3626] = 5'h1b;
assign _c_doomhead[3627] = 5'h17;
assign _c_doomhead[3628] = 5'h17;
assign _c_doomhead[3629] = 5'h1c;
assign _c_doomhead[3630] = 5'h1e;
assign _c_doomhead[3631] = 5'h04;
assign _c_doomhead[3632] = 5'h09;
assign _c_doomhead[3633] = 5'h13;
assign _c_doomhead[3634] = 5'h0f;
assign _c_doomhead[3635] = 5'h0b;
assign _c_doomhead[3636] = 5'h01;
assign _c_doomhead[3637] = 5'h01;
assign _c_doomhead[3638] = 5'h04;
assign _c_doomhead[3639] = 5'h0e;
assign _c_doomhead[3640] = 5'h07;
assign _c_doomhead[3641] = 5'h04;
assign _c_doomhead[3642] = 5'h03;
assign _c_doomhead[3643] = 5'h03;
assign _c_doomhead[3644] = 5'h03;
assign _c_doomhead[3645] = 5'h03;
assign _c_doomhead[3646] = 5'h00;
assign _c_doomhead[3647] = 5'h00;
assign _c_doomhead[3648] = 5'h00;
assign _c_doomhead[3649] = 5'h00;
assign _c_doomhead[3650] = 5'h00;
assign _c_doomhead[3651] = 5'h00;
assign _c_doomhead[3652] = 5'h0b;
assign _c_doomhead[3653] = 5'h1b;
assign _c_doomhead[3654] = 5'h04;
assign _c_doomhead[3655] = 5'h09;
assign _c_doomhead[3656] = 5'h16;
assign _c_doomhead[3657] = 5'h08;
assign _c_doomhead[3658] = 5'h04;
assign _c_doomhead[3659] = 5'h03;
assign _c_doomhead[3660] = 5'h1b;
assign _c_doomhead[3661] = 5'h0c;
assign _c_doomhead[3662] = 5'h04;
assign _c_doomhead[3663] = 5'h04;
assign _c_doomhead[3664] = 5'h0a;
assign _c_doomhead[3665] = 5'h0d;
assign _c_doomhead[3666] = 5'h0c;
assign _c_doomhead[3667] = 5'h09;
assign _c_doomhead[3668] = 5'h08;
assign _c_doomhead[3669] = 5'h08;
assign _c_doomhead[3670] = 5'h0e;
assign _c_doomhead[3671] = 5'h0a;
assign _c_doomhead[3672] = 5'h04;
assign _c_doomhead[3673] = 5'h03;
assign _c_doomhead[3674] = 5'h03;
assign _c_doomhead[3675] = 5'h03;
assign _c_doomhead[3676] = 5'h03;
assign _c_doomhead[3677] = 5'h00;
assign _c_doomhead[3678] = 5'h00;
assign _c_doomhead[3679] = 5'h00;
assign _c_doomhead[3680] = 5'h00;
assign _c_doomhead[3681] = 5'h00;
assign _c_doomhead[3682] = 5'h00;
assign _c_doomhead[3683] = 5'h00;
assign _c_doomhead[3684] = 5'h0b;
assign _c_doomhead[3685] = 5'h18;
assign _c_doomhead[3686] = 5'h01;
assign _c_doomhead[3687] = 5'h0f;
assign _c_doomhead[3688] = 5'h14;
assign _c_doomhead[3689] = 5'h07;
assign _c_doomhead[3690] = 5'h08;
assign _c_doomhead[3691] = 5'h02;
assign _c_doomhead[3692] = 5'h02;
assign _c_doomhead[3693] = 5'h02;
assign _c_doomhead[3694] = 5'h07;
assign _c_doomhead[3695] = 5'h0d;
assign _c_doomhead[3696] = 5'h18;
assign _c_doomhead[3697] = 5'h14;
assign _c_doomhead[3698] = 5'h0f;
assign _c_doomhead[3699] = 5'h08;
assign _c_doomhead[3700] = 5'h01;
assign _c_doomhead[3701] = 5'h08;
assign _c_doomhead[3702] = 5'h01;
assign _c_doomhead[3703] = 5'h04;
assign _c_doomhead[3704] = 5'h0e;
assign _c_doomhead[3705] = 5'h03;
assign _c_doomhead[3706] = 5'h03;
assign _c_doomhead[3707] = 5'h03;
assign _c_doomhead[3708] = 5'h03;
assign _c_doomhead[3709] = 5'h00;
assign _c_doomhead[3710] = 5'h00;
assign _c_doomhead[3711] = 5'h00;
assign _c_doomhead[3712] = 5'h00;
assign _c_doomhead[3713] = 5'h00;
assign _c_doomhead[3714] = 5'h00;
assign _c_doomhead[3715] = 5'h00;
assign _c_doomhead[3716] = 5'h07;
assign _c_doomhead[3717] = 5'h18;
assign _c_doomhead[3718] = 5'h14;
assign _c_doomhead[3719] = 5'h0c;
assign _c_doomhead[3720] = 5'h14;
assign _c_doomhead[3721] = 5'h07;
assign _c_doomhead[3722] = 5'h01;
assign _c_doomhead[3723] = 5'h0d;
assign _c_doomhead[3724] = 5'h1e;
assign _c_doomhead[3725] = 5'h1b;
assign _c_doomhead[3726] = 5'h16;
assign _c_doomhead[3727] = 5'h16;
assign _c_doomhead[3728] = 5'h18;
assign _c_doomhead[3729] = 5'h0c;
assign _c_doomhead[3730] = 5'h09;
assign _c_doomhead[3731] = 5'h08;
assign _c_doomhead[3732] = 5'h09;
assign _c_doomhead[3733] = 5'h08;
assign _c_doomhead[3734] = 5'h01;
assign _c_doomhead[3735] = 5'h15;
assign _c_doomhead[3736] = 5'h15;
assign _c_doomhead[3737] = 5'h03;
assign _c_doomhead[3738] = 5'h03;
assign _c_doomhead[3739] = 5'h03;
assign _c_doomhead[3740] = 5'h03;
assign _c_doomhead[3741] = 5'h00;
assign _c_doomhead[3742] = 5'h00;
assign _c_doomhead[3743] = 5'h00;
assign _c_doomhead[3744] = 5'h00;
assign _c_doomhead[3745] = 5'h00;
assign _c_doomhead[3746] = 5'h00;
assign _c_doomhead[3747] = 5'h00;
assign _c_doomhead[3748] = 5'h08;
assign _c_doomhead[3749] = 5'h0d;
assign _c_doomhead[3750] = 5'h14;
assign _c_doomhead[3751] = 5'h14;
assign _c_doomhead[3752] = 5'h18;
assign _c_doomhead[3753] = 5'h0f;
assign _c_doomhead[3754] = 5'h12;
assign _c_doomhead[3755] = 5'h0b;
assign _c_doomhead[3756] = 5'h09;
assign _c_doomhead[3757] = 5'h1e;
assign _c_doomhead[3758] = 5'h1e;
assign _c_doomhead[3759] = 5'h16;
assign _c_doomhead[3760] = 5'h18;
assign _c_doomhead[3761] = 5'h0a;
assign _c_doomhead[3762] = 5'h08;
assign _c_doomhead[3763] = 5'h08;
assign _c_doomhead[3764] = 5'h0f;
assign _c_doomhead[3765] = 5'h01;
assign _c_doomhead[3766] = 5'h08;
assign _c_doomhead[3767] = 5'h15;
assign _c_doomhead[3768] = 5'h15;
assign _c_doomhead[3769] = 5'h03;
assign _c_doomhead[3770] = 5'h03;
assign _c_doomhead[3771] = 5'h03;
assign _c_doomhead[3772] = 5'h03;
assign _c_doomhead[3773] = 5'h00;
assign _c_doomhead[3774] = 5'h00;
assign _c_doomhead[3775] = 5'h00;
assign _c_doomhead[3776] = 5'h00;
assign _c_doomhead[3777] = 5'h00;
assign _c_doomhead[3778] = 5'h00;
assign _c_doomhead[3779] = 5'h00;
assign _c_doomhead[3780] = 5'h00;
assign _c_doomhead[3781] = 5'h01;
assign _c_doomhead[3782] = 5'h0d;
assign _c_doomhead[3783] = 5'h0f;
assign _c_doomhead[3784] = 5'h18;
assign _c_doomhead[3785] = 5'h0a;
assign _c_doomhead[3786] = 5'h06;
assign _c_doomhead[3787] = 5'h04;
assign _c_doomhead[3788] = 5'h08;
assign _c_doomhead[3789] = 5'h03;
assign _c_doomhead[3790] = 5'h1e;
assign _c_doomhead[3791] = 5'h19;
assign _c_doomhead[3792] = 5'h12;
assign _c_doomhead[3793] = 5'h0f;
assign _c_doomhead[3794] = 5'h08;
assign _c_doomhead[3795] = 5'h08;
assign _c_doomhead[3796] = 5'h0f;
assign _c_doomhead[3797] = 5'h09;
assign _c_doomhead[3798] = 5'h07;
assign _c_doomhead[3799] = 5'h15;
assign _c_doomhead[3800] = 5'h01;
assign _c_doomhead[3801] = 5'h03;
assign _c_doomhead[3802] = 5'h03;
assign _c_doomhead[3803] = 5'h03;
assign _c_doomhead[3804] = 5'h00;
assign _c_doomhead[3805] = 5'h00;
assign _c_doomhead[3806] = 5'h00;
assign _c_doomhead[3807] = 5'h00;
assign _c_doomhead[3808] = 5'h00;
assign _c_doomhead[3809] = 5'h00;
assign _c_doomhead[3810] = 5'h00;
assign _c_doomhead[3811] = 5'h00;
assign _c_doomhead[3812] = 5'h00;
assign _c_doomhead[3813] = 5'h04;
assign _c_doomhead[3814] = 5'h0b;
assign _c_doomhead[3815] = 5'h01;
assign _c_doomhead[3816] = 5'h0a;
assign _c_doomhead[3817] = 5'h04;
assign _c_doomhead[3818] = 5'h1c;
assign _c_doomhead[3819] = 5'h1c;
assign _c_doomhead[3820] = 5'h09;
assign _c_doomhead[3821] = 5'h1a;
assign _c_doomhead[3822] = 5'h03;
assign _c_doomhead[3823] = 5'h0c;
assign _c_doomhead[3824] = 5'h0d;
assign _c_doomhead[3825] = 5'h0c;
assign _c_doomhead[3826] = 5'h08;
assign _c_doomhead[3827] = 5'h01;
assign _c_doomhead[3828] = 5'h0b;
assign _c_doomhead[3829] = 5'h07;
assign _c_doomhead[3830] = 5'h07;
assign _c_doomhead[3831] = 5'h01;
assign _c_doomhead[3832] = 5'h01;
assign _c_doomhead[3833] = 5'h15;
assign _c_doomhead[3834] = 5'h03;
assign _c_doomhead[3835] = 5'h03;
assign _c_doomhead[3836] = 5'h00;
assign _c_doomhead[3837] = 5'h00;
assign _c_doomhead[3838] = 5'h00;
assign _c_doomhead[3839] = 5'h00;
assign _c_doomhead[3840] = 5'h00;
assign _c_doomhead[3841] = 5'h00;
assign _c_doomhead[3842] = 5'h00;
assign _c_doomhead[3843] = 5'h00;
assign _c_doomhead[3844] = 5'h00;
assign _c_doomhead[3845] = 5'h00;
assign _c_doomhead[3846] = 5'h07;
assign _c_doomhead[3847] = 5'h1a;
assign _c_doomhead[3848] = 5'h1c;
assign _c_doomhead[3849] = 5'h03;
assign _c_doomhead[3850] = 5'h1c;
assign _c_doomhead[3851] = 5'h1c;
assign _c_doomhead[3852] = 5'h0c;
assign _c_doomhead[3853] = 5'h14;
assign _c_doomhead[3854] = 5'h1a;
assign _c_doomhead[3855] = 5'h1e;
assign _c_doomhead[3856] = 5'h0c;
assign _c_doomhead[3857] = 5'h0c;
assign _c_doomhead[3858] = 5'h01;
assign _c_doomhead[3859] = 5'h07;
assign _c_doomhead[3860] = 5'h07;
assign _c_doomhead[3861] = 5'h07;
assign _c_doomhead[3862] = 5'h15;
assign _c_doomhead[3863] = 5'h01;
assign _c_doomhead[3864] = 5'h07;
assign _c_doomhead[3865] = 5'h15;
assign _c_doomhead[3866] = 5'h00;
assign _c_doomhead[3867] = 5'h00;
assign _c_doomhead[3868] = 5'h00;
assign _c_doomhead[3869] = 5'h00;
assign _c_doomhead[3870] = 5'h00;
assign _c_doomhead[3871] = 5'h00;
assign _c_doomhead[3872] = 5'h00;
assign _c_doomhead[3873] = 5'h00;
assign _c_doomhead[3874] = 5'h00;
assign _c_doomhead[3875] = 5'h00;
assign _c_doomhead[3876] = 5'h00;
assign _c_doomhead[3877] = 5'h00;
assign _c_doomhead[3878] = 5'h01;
assign _c_doomhead[3879] = 5'h1d;
assign _c_doomhead[3880] = 5'h1c;
assign _c_doomhead[3881] = 5'h1d;
assign _c_doomhead[3882] = 5'h1e;
assign _c_doomhead[3883] = 5'h1e;
assign _c_doomhead[3884] = 5'h19;
assign _c_doomhead[3885] = 5'h0c;
assign _c_doomhead[3886] = 5'h1e;
assign _c_doomhead[3887] = 5'h1a;
assign _c_doomhead[3888] = 5'h0c;
assign _c_doomhead[3889] = 5'h0f;
assign _c_doomhead[3890] = 5'h01;
assign _c_doomhead[3891] = 5'h07;
assign _c_doomhead[3892] = 5'h07;
assign _c_doomhead[3893] = 5'h08;
assign _c_doomhead[3894] = 5'h02;
assign _c_doomhead[3895] = 5'h01;
assign _c_doomhead[3896] = 5'h00;
assign _c_doomhead[3897] = 5'h00;
assign _c_doomhead[3898] = 5'h00;
assign _c_doomhead[3899] = 5'h00;
assign _c_doomhead[3900] = 5'h00;
assign _c_doomhead[3901] = 5'h00;
assign _c_doomhead[3902] = 5'h00;
assign _c_doomhead[3903] = 5'h00;
assign _c_doomhead[3904] = 5'h00;
assign _c_doomhead[3905] = 5'h00;
assign _c_doomhead[3906] = 5'h00;
assign _c_doomhead[3907] = 5'h00;
assign _c_doomhead[3908] = 5'h00;
assign _c_doomhead[3909] = 5'h00;
assign _c_doomhead[3910] = 5'h04;
assign _c_doomhead[3911] = 5'h1e;
assign _c_doomhead[3912] = 5'h1c;
assign _c_doomhead[3913] = 5'h1c;
assign _c_doomhead[3914] = 5'h1a;
assign _c_doomhead[3915] = 5'h1b;
assign _c_doomhead[3916] = 5'h1c;
assign _c_doomhead[3917] = 5'h1c;
assign _c_doomhead[3918] = 5'h1d;
assign _c_doomhead[3919] = 5'h1a;
assign _c_doomhead[3920] = 5'h1e;
assign _c_doomhead[3921] = 5'h0f;
assign _c_doomhead[3922] = 5'h09;
assign _c_doomhead[3923] = 5'h07;
assign _c_doomhead[3924] = 5'h15;
assign _c_doomhead[3925] = 5'h02;
assign _c_doomhead[3926] = 5'h04;
assign _c_doomhead[3927] = 5'h00;
assign _c_doomhead[3928] = 5'h00;
assign _c_doomhead[3929] = 5'h00;
assign _c_doomhead[3930] = 5'h00;
assign _c_doomhead[3931] = 5'h00;
assign _c_doomhead[3932] = 5'h00;
assign _c_doomhead[3933] = 5'h00;
assign _c_doomhead[3934] = 5'h00;
assign _c_doomhead[3935] = 5'h00;
assign _c_doomhead[3936] = 5'h00;
assign _c_doomhead[3937] = 5'h00;
assign _c_doomhead[3938] = 5'h00;
assign _c_doomhead[3939] = 5'h00;
assign _c_doomhead[3940] = 5'h00;
assign _c_doomhead[3941] = 5'h00;
assign _c_doomhead[3942] = 5'h00;
assign _c_doomhead[3943] = 5'h01;
assign _c_doomhead[3944] = 5'h1a;
assign _c_doomhead[3945] = 5'h1e;
assign _c_doomhead[3946] = 5'h1e;
assign _c_doomhead[3947] = 5'h1d;
assign _c_doomhead[3948] = 5'h0c;
assign _c_doomhead[3949] = 5'h0b;
assign _c_doomhead[3950] = 5'h1e;
assign _c_doomhead[3951] = 5'h1b;
assign _c_doomhead[3952] = 5'h1d;
assign _c_doomhead[3953] = 5'h0f;
assign _c_doomhead[3954] = 5'h09;
assign _c_doomhead[3955] = 5'h07;
assign _c_doomhead[3956] = 5'h15;
assign _c_doomhead[3957] = 5'h04;
assign _c_doomhead[3958] = 5'h00;
assign _c_doomhead[3959] = 5'h00;
assign _c_doomhead[3960] = 5'h00;
assign _c_doomhead[3961] = 5'h00;
assign _c_doomhead[3962] = 5'h00;
assign _c_doomhead[3963] = 5'h00;
assign _c_doomhead[3964] = 5'h00;
assign _c_doomhead[3965] = 5'h00;
assign _c_doomhead[3966] = 5'h00;
assign _c_doomhead[3967] = 5'h00;
assign _c_doomhead[3968] = 5'h00;
assign _c_doomhead[3969] = 5'h00;
assign _c_doomhead[3970] = 5'h00;
assign _c_doomhead[3971] = 5'h00;
assign _c_doomhead[3972] = 5'h00;
assign _c_doomhead[3973] = 5'h00;
assign _c_doomhead[3974] = 5'h00;
assign _c_doomhead[3975] = 5'h01;
assign _c_doomhead[3976] = 5'h09;
assign _c_doomhead[3977] = 5'h1c;
assign _c_doomhead[3978] = 5'h1c;
assign _c_doomhead[3979] = 5'h1a;
assign _c_doomhead[3980] = 5'h1a;
assign _c_doomhead[3981] = 5'h07;
assign _c_doomhead[3982] = 5'h0b;
assign _c_doomhead[3983] = 5'h1b;
assign _c_doomhead[3984] = 5'h1d;
assign _c_doomhead[3985] = 5'h0b;
assign _c_doomhead[3986] = 5'h07;
assign _c_doomhead[3987] = 5'h02;
assign _c_doomhead[3988] = 5'h05;
assign _c_doomhead[3989] = 5'h00;
assign _c_doomhead[3990] = 5'h00;
assign _c_doomhead[3991] = 5'h00;
assign _c_doomhead[3992] = 5'h00;
assign _c_doomhead[3993] = 5'h00;
assign _c_doomhead[3994] = 5'h00;
assign _c_doomhead[3995] = 5'h00;
assign _c_doomhead[3996] = 5'h00;
assign _c_doomhead[3997] = 5'h00;
assign _c_doomhead[3998] = 5'h00;
assign _c_doomhead[3999] = 5'h00;
assign _c_doomhead[4000] = 5'h00;
assign _c_doomhead[4001] = 5'h00;
assign _c_doomhead[4002] = 5'h00;
assign _c_doomhead[4003] = 5'h00;
assign _c_doomhead[4004] = 5'h00;
assign _c_doomhead[4005] = 5'h00;
assign _c_doomhead[4006] = 5'h00;
assign _c_doomhead[4007] = 5'h04;
assign _c_doomhead[4008] = 5'h01;
assign _c_doomhead[4009] = 5'h1a;
assign _c_doomhead[4010] = 5'h1e;
assign _c_doomhead[4011] = 5'h1a;
assign _c_doomhead[4012] = 5'h1d;
assign _c_doomhead[4013] = 5'h0f;
assign _c_doomhead[4014] = 5'h0f;
assign _c_doomhead[4015] = 5'h1b;
assign _c_doomhead[4016] = 5'h1c;
assign _c_doomhead[4017] = 5'h15;
assign _c_doomhead[4018] = 5'h05;
assign _c_doomhead[4019] = 5'h05;
assign _c_doomhead[4020] = 5'h00;
assign _c_doomhead[4021] = 5'h00;
assign _c_doomhead[4022] = 5'h00;
assign _c_doomhead[4023] = 5'h00;
assign _c_doomhead[4024] = 5'h00;
assign _c_doomhead[4025] = 5'h00;
assign _c_doomhead[4026] = 5'h00;
assign _c_doomhead[4027] = 5'h00;
assign _c_doomhead[4028] = 5'h00;
assign _c_doomhead[4029] = 5'h00;
assign _c_doomhead[4030] = 5'h00;
assign _c_doomhead[4031] = 5'h00;
assign _c_doomhead[4032] = 5'h00;
assign _c_doomhead[4033] = 5'h00;
assign _c_doomhead[4034] = 5'h00;
assign _c_doomhead[4035] = 5'h00;
assign _c_doomhead[4036] = 5'h00;
assign _c_doomhead[4037] = 5'h00;
assign _c_doomhead[4038] = 5'h00;
assign _c_doomhead[4039] = 5'h00;
assign _c_doomhead[4040] = 5'h04;
assign _c_doomhead[4041] = 5'h1a;
assign _c_doomhead[4042] = 5'h1c;
assign _c_doomhead[4043] = 5'h1c;
assign _c_doomhead[4044] = 5'h1d;
assign _c_doomhead[4045] = 5'h09;
assign _c_doomhead[4046] = 5'h01;
assign _c_doomhead[4047] = 5'h1b;
assign _c_doomhead[4048] = 5'h1c;
assign _c_doomhead[4049] = 5'h05;
assign _c_doomhead[4050] = 5'h05;
assign _c_doomhead[4051] = 5'h00;
assign _c_doomhead[4052] = 5'h00;
assign _c_doomhead[4053] = 5'h00;
assign _c_doomhead[4054] = 5'h00;
assign _c_doomhead[4055] = 5'h00;
assign _c_doomhead[4056] = 5'h00;
assign _c_doomhead[4057] = 5'h00;
assign _c_doomhead[4058] = 5'h00;
assign _c_doomhead[4059] = 5'h00;
assign _c_doomhead[4060] = 5'h00;
assign _c_doomhead[4061] = 5'h00;
assign _c_doomhead[4062] = 5'h00;
assign _c_doomhead[4063] = 5'h00;
assign _c_doomhead[4064] = 5'h00;
assign _c_doomhead[4065] = 5'h00;
assign _c_doomhead[4066] = 5'h00;
assign _c_doomhead[4067] = 5'h00;
assign _c_doomhead[4068] = 5'h00;
assign _c_doomhead[4069] = 5'h00;
assign _c_doomhead[4070] = 5'h00;
assign _c_doomhead[4071] = 5'h00;
assign _c_doomhead[4072] = 5'h00;
assign _c_doomhead[4073] = 5'h00;
assign _c_doomhead[4074] = 5'h00;
assign _c_doomhead[4075] = 5'h00;
assign _c_doomhead[4076] = 5'h00;
assign _c_doomhead[4077] = 5'h00;
assign _c_doomhead[4078] = 5'h00;
assign _c_doomhead[4079] = 5'h00;
assign _c_doomhead[4080] = 5'h00;
assign _c_doomhead[4081] = 5'h00;
assign _c_doomhead[4082] = 5'h00;
assign _c_doomhead[4083] = 5'h00;
assign _c_doomhead[4084] = 5'h00;
assign _c_doomhead[4085] = 5'h00;
assign _c_doomhead[4086] = 5'h00;
assign _c_doomhead[4087] = 5'h00;
assign _c_doomhead[4088] = 5'h00;
assign _c_doomhead[4089] = 5'h00;
assign _c_doomhead[4090] = 5'h00;
assign _c_doomhead[4091] = 5'h00;
assign _c_doomhead[4092] = 5'h00;
assign _c_doomhead[4093] = 5'h00;
assign _c_doomhead[4094] = 5'h00;
assign _c_doomhead[4095] = 5'h00;
assign _c_doomhead[4096] = 5'h00;
assign _c_doomhead[4097] = 5'h00;
assign _c_doomhead[4098] = 5'h00;
assign _c_doomhead[4099] = 5'h00;
assign _c_doomhead[4100] = 5'h00;
assign _c_doomhead[4101] = 5'h00;
assign _c_doomhead[4102] = 5'h00;
assign _c_doomhead[4103] = 5'h00;
assign _c_doomhead[4104] = 5'h00;
assign _c_doomhead[4105] = 5'h02;
assign _c_doomhead[4106] = 5'h04;
assign _c_doomhead[4107] = 5'h04;
assign _c_doomhead[4108] = 5'h06;
assign _c_doomhead[4109] = 5'h06;
assign _c_doomhead[4110] = 5'h08;
assign _c_doomhead[4111] = 5'h08;
assign _c_doomhead[4112] = 5'h08;
assign _c_doomhead[4113] = 5'h04;
assign _c_doomhead[4114] = 5'h02;
assign _c_doomhead[4115] = 5'h02;
assign _c_doomhead[4116] = 5'h00;
assign _c_doomhead[4117] = 5'h00;
assign _c_doomhead[4118] = 5'h00;
assign _c_doomhead[4119] = 5'h00;
assign _c_doomhead[4120] = 5'h00;
assign _c_doomhead[4121] = 5'h00;
assign _c_doomhead[4122] = 5'h00;
assign _c_doomhead[4123] = 5'h00;
assign _c_doomhead[4124] = 5'h00;
assign _c_doomhead[4125] = 5'h00;
assign _c_doomhead[4126] = 5'h00;
assign _c_doomhead[4127] = 5'h00;
assign _c_doomhead[4128] = 5'h00;
assign _c_doomhead[4129] = 5'h00;
assign _c_doomhead[4130] = 5'h00;
assign _c_doomhead[4131] = 5'h00;
assign _c_doomhead[4132] = 5'h00;
assign _c_doomhead[4133] = 5'h00;
assign _c_doomhead[4134] = 5'h00;
assign _c_doomhead[4135] = 5'h05;
assign _c_doomhead[4136] = 5'h05;
assign _c_doomhead[4137] = 5'h02;
assign _c_doomhead[4138] = 5'h04;
assign _c_doomhead[4139] = 5'h06;
assign _c_doomhead[4140] = 5'h08;
assign _c_doomhead[4141] = 5'h01;
assign _c_doomhead[4142] = 5'h07;
assign _c_doomhead[4143] = 5'h07;
assign _c_doomhead[4144] = 5'h0a;
assign _c_doomhead[4145] = 5'h0a;
assign _c_doomhead[4146] = 5'h01;
assign _c_doomhead[4147] = 5'h08;
assign _c_doomhead[4148] = 5'h04;
assign _c_doomhead[4149] = 5'h02;
assign _c_doomhead[4150] = 5'h00;
assign _c_doomhead[4151] = 5'h00;
assign _c_doomhead[4152] = 5'h00;
assign _c_doomhead[4153] = 5'h00;
assign _c_doomhead[4154] = 5'h00;
assign _c_doomhead[4155] = 5'h00;
assign _c_doomhead[4156] = 5'h00;
assign _c_doomhead[4157] = 5'h00;
assign _c_doomhead[4158] = 5'h00;
assign _c_doomhead[4159] = 5'h00;
assign _c_doomhead[4160] = 5'h00;
assign _c_doomhead[4161] = 5'h00;
assign _c_doomhead[4162] = 5'h00;
assign _c_doomhead[4163] = 5'h00;
assign _c_doomhead[4164] = 5'h00;
assign _c_doomhead[4165] = 5'h10;
assign _c_doomhead[4166] = 5'h10;
assign _c_doomhead[4167] = 5'h05;
assign _c_doomhead[4168] = 5'h05;
assign _c_doomhead[4169] = 5'h02;
assign _c_doomhead[4170] = 5'h02;
assign _c_doomhead[4171] = 5'h06;
assign _c_doomhead[4172] = 5'h08;
assign _c_doomhead[4173] = 5'h01;
assign _c_doomhead[4174] = 5'h07;
assign _c_doomhead[4175] = 5'h07;
assign _c_doomhead[4176] = 5'h07;
assign _c_doomhead[4177] = 5'h07;
assign _c_doomhead[4178] = 5'h01;
assign _c_doomhead[4179] = 5'h08;
assign _c_doomhead[4180] = 5'h04;
assign _c_doomhead[4181] = 5'h02;
assign _c_doomhead[4182] = 5'h05;
assign _c_doomhead[4183] = 5'h03;
assign _c_doomhead[4184] = 5'h00;
assign _c_doomhead[4185] = 5'h00;
assign _c_doomhead[4186] = 5'h00;
assign _c_doomhead[4187] = 5'h00;
assign _c_doomhead[4188] = 5'h00;
assign _c_doomhead[4189] = 5'h00;
assign _c_doomhead[4190] = 5'h00;
assign _c_doomhead[4191] = 5'h00;
assign _c_doomhead[4192] = 5'h00;
assign _c_doomhead[4193] = 5'h00;
assign _c_doomhead[4194] = 5'h00;
assign _c_doomhead[4195] = 5'h00;
assign _c_doomhead[4196] = 5'h10;
assign _c_doomhead[4197] = 5'h03;
assign _c_doomhead[4198] = 5'h05;
assign _c_doomhead[4199] = 5'h10;
assign _c_doomhead[4200] = 5'h05;
assign _c_doomhead[4201] = 5'h05;
assign _c_doomhead[4202] = 5'h02;
assign _c_doomhead[4203] = 5'h02;
assign _c_doomhead[4204] = 5'h02;
assign _c_doomhead[4205] = 5'h06;
assign _c_doomhead[4206] = 5'h08;
assign _c_doomhead[4207] = 5'h01;
assign _c_doomhead[4208] = 5'h07;
assign _c_doomhead[4209] = 5'h0a;
assign _c_doomhead[4210] = 5'h0f;
assign _c_doomhead[4211] = 5'h0f;
assign _c_doomhead[4212] = 5'h0a;
assign _c_doomhead[4213] = 5'h01;
assign _c_doomhead[4214] = 5'h02;
assign _c_doomhead[4215] = 5'h05;
assign _c_doomhead[4216] = 5'h05;
assign _c_doomhead[4217] = 5'h00;
assign _c_doomhead[4218] = 5'h00;
assign _c_doomhead[4219] = 5'h00;
assign _c_doomhead[4220] = 5'h00;
assign _c_doomhead[4221] = 5'h00;
assign _c_doomhead[4222] = 5'h00;
assign _c_doomhead[4223] = 5'h00;
assign _c_doomhead[4224] = 5'h00;
assign _c_doomhead[4225] = 5'h00;
assign _c_doomhead[4226] = 5'h00;
assign _c_doomhead[4227] = 5'h03;
assign _c_doomhead[4228] = 5'h10;
assign _c_doomhead[4229] = 5'h05;
assign _c_doomhead[4230] = 5'h10;
assign _c_doomhead[4231] = 5'h10;
assign _c_doomhead[4232] = 5'h05;
assign _c_doomhead[4233] = 5'h05;
assign _c_doomhead[4234] = 5'h02;
assign _c_doomhead[4235] = 5'h02;
assign _c_doomhead[4236] = 5'h02;
assign _c_doomhead[4237] = 5'h02;
assign _c_doomhead[4238] = 5'h06;
assign _c_doomhead[4239] = 5'h08;
assign _c_doomhead[4240] = 5'h01;
assign _c_doomhead[4241] = 5'h07;
assign _c_doomhead[4242] = 5'h07;
assign _c_doomhead[4243] = 5'h07;
assign _c_doomhead[4244] = 5'h07;
assign _c_doomhead[4245] = 5'h07;
assign _c_doomhead[4246] = 5'h01;
assign _c_doomhead[4247] = 5'h02;
assign _c_doomhead[4248] = 5'h05;
assign _c_doomhead[4249] = 5'h05;
assign _c_doomhead[4250] = 5'h00;
assign _c_doomhead[4251] = 5'h00;
assign _c_doomhead[4252] = 5'h00;
assign _c_doomhead[4253] = 5'h00;
assign _c_doomhead[4254] = 5'h00;
assign _c_doomhead[4255] = 5'h00;
assign _c_doomhead[4256] = 5'h00;
assign _c_doomhead[4257] = 5'h00;
assign _c_doomhead[4258] = 5'h00;
assign _c_doomhead[4259] = 5'h10;
assign _c_doomhead[4260] = 5'h10;
assign _c_doomhead[4261] = 5'h10;
assign _c_doomhead[4262] = 5'h10;
assign _c_doomhead[4263] = 5'h05;
assign _c_doomhead[4264] = 5'h05;
assign _c_doomhead[4265] = 5'h05;
assign _c_doomhead[4266] = 5'h05;
assign _c_doomhead[4267] = 5'h02;
assign _c_doomhead[4268] = 5'h02;
assign _c_doomhead[4269] = 5'h02;
assign _c_doomhead[4270] = 5'h04;
assign _c_doomhead[4271] = 5'h06;
assign _c_doomhead[4272] = 5'h06;
assign _c_doomhead[4273] = 5'h01;
assign _c_doomhead[4274] = 5'h01;
assign _c_doomhead[4275] = 5'h06;
assign _c_doomhead[4276] = 5'h06;
assign _c_doomhead[4277] = 5'h06;
assign _c_doomhead[4278] = 5'h06;
assign _c_doomhead[4279] = 5'h04;
assign _c_doomhead[4280] = 5'h06;
assign _c_doomhead[4281] = 5'h06;
assign _c_doomhead[4282] = 5'h02;
assign _c_doomhead[4283] = 5'h00;
assign _c_doomhead[4284] = 5'h00;
assign _c_doomhead[4285] = 5'h00;
assign _c_doomhead[4286] = 5'h00;
assign _c_doomhead[4287] = 5'h00;
assign _c_doomhead[4288] = 5'h00;
assign _c_doomhead[4289] = 5'h00;
assign _c_doomhead[4290] = 5'h03;
assign _c_doomhead[4291] = 5'h10;
assign _c_doomhead[4292] = 5'h10;
assign _c_doomhead[4293] = 5'h10;
assign _c_doomhead[4294] = 5'h05;
assign _c_doomhead[4295] = 5'h05;
assign _c_doomhead[4296] = 5'h10;
assign _c_doomhead[4297] = 5'h10;
assign _c_doomhead[4298] = 5'h0e;
assign _c_doomhead[4299] = 5'h04;
assign _c_doomhead[4300] = 5'h0e;
assign _c_doomhead[4301] = 5'h0e;
assign _c_doomhead[4302] = 5'h02;
assign _c_doomhead[4303] = 5'h09;
assign _c_doomhead[4304] = 5'h01;
assign _c_doomhead[4305] = 5'h04;
assign _c_doomhead[4306] = 5'h04;
assign _c_doomhead[4307] = 5'h04;
assign _c_doomhead[4308] = 5'h06;
assign _c_doomhead[4309] = 5'h01;
assign _c_doomhead[4310] = 5'h01;
assign _c_doomhead[4311] = 5'h08;
assign _c_doomhead[4312] = 5'h08;
assign _c_doomhead[4313] = 5'h07;
assign _c_doomhead[4314] = 5'h08;
assign _c_doomhead[4315] = 5'h04;
assign _c_doomhead[4316] = 5'h00;
assign _c_doomhead[4317] = 5'h00;
assign _c_doomhead[4318] = 5'h00;
assign _c_doomhead[4319] = 5'h00;
assign _c_doomhead[4320] = 5'h00;
assign _c_doomhead[4321] = 5'h00;
assign _c_doomhead[4322] = 5'h03;
assign _c_doomhead[4323] = 5'h03;
assign _c_doomhead[4324] = 5'h03;
assign _c_doomhead[4325] = 5'h05;
assign _c_doomhead[4326] = 5'h03;
assign _c_doomhead[4327] = 5'h10;
assign _c_doomhead[4328] = 5'h05;
assign _c_doomhead[4329] = 5'h04;
assign _c_doomhead[4330] = 5'h04;
assign _c_doomhead[4331] = 5'h0e;
assign _c_doomhead[4332] = 5'h04;
assign _c_doomhead[4333] = 5'h01;
assign _c_doomhead[4334] = 5'h15;
assign _c_doomhead[4335] = 5'h02;
assign _c_doomhead[4336] = 5'h02;
assign _c_doomhead[4337] = 5'h05;
assign _c_doomhead[4338] = 5'h05;
assign _c_doomhead[4339] = 5'h06;
assign _c_doomhead[4340] = 5'h04;
assign _c_doomhead[4341] = 5'h02;
assign _c_doomhead[4342] = 5'h04;
assign _c_doomhead[4343] = 5'h08;
assign _c_doomhead[4344] = 5'h07;
assign _c_doomhead[4345] = 5'h10;
assign _c_doomhead[4346] = 5'h10;
assign _c_doomhead[4347] = 5'h10;
assign _c_doomhead[4348] = 5'h11;
assign _c_doomhead[4349] = 5'h00;
assign _c_doomhead[4350] = 5'h00;
assign _c_doomhead[4351] = 5'h00;
assign _c_doomhead[4352] = 5'h00;
assign _c_doomhead[4353] = 5'h03;
assign _c_doomhead[4354] = 5'h03;
assign _c_doomhead[4355] = 5'h03;
assign _c_doomhead[4356] = 5'h03;
assign _c_doomhead[4357] = 5'h03;
assign _c_doomhead[4358] = 5'h10;
assign _c_doomhead[4359] = 5'h05;
assign _c_doomhead[4360] = 5'h04;
assign _c_doomhead[4361] = 5'h05;
assign _c_doomhead[4362] = 5'h02;
assign _c_doomhead[4363] = 5'h01;
assign _c_doomhead[4364] = 5'h04;
assign _c_doomhead[4365] = 5'h10;
assign _c_doomhead[4366] = 5'h10;
assign _c_doomhead[4367] = 5'h03;
assign _c_doomhead[4368] = 5'h10;
assign _c_doomhead[4369] = 5'h05;
assign _c_doomhead[4370] = 5'h04;
assign _c_doomhead[4371] = 5'h05;
assign _c_doomhead[4372] = 5'h04;
assign _c_doomhead[4373] = 5'h04;
assign _c_doomhead[4374] = 5'h07;
assign _c_doomhead[4375] = 5'h04;
assign _c_doomhead[4376] = 5'h02;
assign _c_doomhead[4377] = 5'h11;
assign _c_doomhead[4378] = 5'h11;
assign _c_doomhead[4379] = 5'h11;
assign _c_doomhead[4380] = 5'h05;
assign _c_doomhead[4381] = 5'h00;
assign _c_doomhead[4382] = 5'h00;
assign _c_doomhead[4383] = 5'h00;
assign _c_doomhead[4384] = 5'h00;
assign _c_doomhead[4385] = 5'h03;
assign _c_doomhead[4386] = 5'h03;
assign _c_doomhead[4387] = 5'h03;
assign _c_doomhead[4388] = 5'h03;
assign _c_doomhead[4389] = 5'h03;
assign _c_doomhead[4390] = 5'h03;
assign _c_doomhead[4391] = 5'h03;
assign _c_doomhead[4392] = 5'h03;
assign _c_doomhead[4393] = 5'h03;
assign _c_doomhead[4394] = 5'h03;
assign _c_doomhead[4395] = 5'h02;
assign _c_doomhead[4396] = 5'h02;
assign _c_doomhead[4397] = 5'h08;
assign _c_doomhead[4398] = 5'h07;
assign _c_doomhead[4399] = 5'h09;
assign _c_doomhead[4400] = 5'h0a;
assign _c_doomhead[4401] = 5'h1c;
assign _c_doomhead[4402] = 5'h1a;
assign _c_doomhead[4403] = 5'h1c;
assign _c_doomhead[4404] = 5'h10;
assign _c_doomhead[4405] = 5'h04;
assign _c_doomhead[4406] = 5'h04;
assign _c_doomhead[4407] = 5'h11;
assign _c_doomhead[4408] = 5'h02;
assign _c_doomhead[4409] = 5'h05;
assign _c_doomhead[4410] = 5'h03;
assign _c_doomhead[4411] = 5'h11;
assign _c_doomhead[4412] = 5'h00;
assign _c_doomhead[4413] = 5'h00;
assign _c_doomhead[4414] = 5'h00;
assign _c_doomhead[4415] = 5'h00;
assign _c_doomhead[4416] = 5'h00;
assign _c_doomhead[4417] = 5'h03;
assign _c_doomhead[4418] = 5'h03;
assign _c_doomhead[4419] = 5'h03;
assign _c_doomhead[4420] = 5'h03;
assign _c_doomhead[4421] = 5'h03;
assign _c_doomhead[4422] = 5'h03;
assign _c_doomhead[4423] = 5'h03;
assign _c_doomhead[4424] = 5'h03;
assign _c_doomhead[4425] = 5'h03;
assign _c_doomhead[4426] = 5'h05;
assign _c_doomhead[4427] = 5'h02;
assign _c_doomhead[4428] = 5'h01;
assign _c_doomhead[4429] = 5'h0b;
assign _c_doomhead[4430] = 5'h0b;
assign _c_doomhead[4431] = 5'h0f;
assign _c_doomhead[4432] = 5'h14;
assign _c_doomhead[4433] = 5'h1b;
assign _c_doomhead[4434] = 5'h1d;
assign _c_doomhead[4435] = 5'h1b;
assign _c_doomhead[4436] = 5'h1c;
assign _c_doomhead[4437] = 5'h02;
assign _c_doomhead[4438] = 5'h0b;
assign _c_doomhead[4439] = 5'h14;
assign _c_doomhead[4440] = 5'h05;
assign _c_doomhead[4441] = 5'h1c;
assign _c_doomhead[4442] = 5'h05;
assign _c_doomhead[4443] = 5'h05;
assign _c_doomhead[4444] = 5'h00;
assign _c_doomhead[4445] = 5'h00;
assign _c_doomhead[4446] = 5'h00;
assign _c_doomhead[4447] = 5'h00;
assign _c_doomhead[4448] = 5'h00;
assign _c_doomhead[4449] = 5'h03;
assign _c_doomhead[4450] = 5'h03;
assign _c_doomhead[4451] = 5'h03;
assign _c_doomhead[4452] = 5'h03;
assign _c_doomhead[4453] = 5'h03;
assign _c_doomhead[4454] = 5'h03;
assign _c_doomhead[4455] = 5'h03;
assign _c_doomhead[4456] = 5'h03;
assign _c_doomhead[4457] = 5'h05;
assign _c_doomhead[4458] = 5'h02;
assign _c_doomhead[4459] = 5'h02;
assign _c_doomhead[4460] = 5'h01;
assign _c_doomhead[4461] = 5'h0b;
assign _c_doomhead[4462] = 5'h0f;
assign _c_doomhead[4463] = 5'h0d;
assign _c_doomhead[4464] = 5'h19;
assign _c_doomhead[4465] = 5'h1b;
assign _c_doomhead[4466] = 5'h1b;
assign _c_doomhead[4467] = 5'h1c;
assign _c_doomhead[4468] = 5'h0d;
assign _c_doomhead[4469] = 5'h0d;
assign _c_doomhead[4470] = 5'h09;
assign _c_doomhead[4471] = 5'h0d;
assign _c_doomhead[4472] = 5'h1e;
assign _c_doomhead[4473] = 5'h10;
assign _c_doomhead[4474] = 5'h05;
assign _c_doomhead[4475] = 5'h00;
assign _c_doomhead[4476] = 5'h00;
assign _c_doomhead[4477] = 5'h00;
assign _c_doomhead[4478] = 5'h00;
assign _c_doomhead[4479] = 5'h00;
assign _c_doomhead[4480] = 5'h00;
assign _c_doomhead[4481] = 5'h03;
assign _c_doomhead[4482] = 5'h03;
assign _c_doomhead[4483] = 5'h03;
assign _c_doomhead[4484] = 5'h03;
assign _c_doomhead[4485] = 5'h04;
assign _c_doomhead[4486] = 5'h04;
assign _c_doomhead[4487] = 5'h04;
assign _c_doomhead[4488] = 5'h04;
assign _c_doomhead[4489] = 5'h05;
assign _c_doomhead[4490] = 5'h05;
assign _c_doomhead[4491] = 5'h02;
assign _c_doomhead[4492] = 5'h01;
assign _c_doomhead[4493] = 5'h0b;
assign _c_doomhead[4494] = 5'h0a;
assign _c_doomhead[4495] = 5'h0d;
assign _c_doomhead[4496] = 5'h0d;
assign _c_doomhead[4497] = 5'h1b;
assign _c_doomhead[4498] = 5'h1e;
assign _c_doomhead[4499] = 5'h0d;
assign _c_doomhead[4500] = 5'h0d;
assign _c_doomhead[4501] = 5'h0d;
assign _c_doomhead[4502] = 5'h0d;
assign _c_doomhead[4503] = 5'h0b;
assign _c_doomhead[4504] = 5'h1e;
assign _c_doomhead[4505] = 5'h1c;
assign _c_doomhead[4506] = 5'h09;
assign _c_doomhead[4507] = 5'h00;
assign _c_doomhead[4508] = 5'h00;
assign _c_doomhead[4509] = 5'h00;
assign _c_doomhead[4510] = 5'h00;
assign _c_doomhead[4511] = 5'h00;
assign _c_doomhead[4512] = 5'h00;
assign _c_doomhead[4513] = 5'h03;
assign _c_doomhead[4514] = 5'h03;
assign _c_doomhead[4515] = 5'h03;
assign _c_doomhead[4516] = 5'h08;
assign _c_doomhead[4517] = 5'h08;
assign _c_doomhead[4518] = 5'h07;
assign _c_doomhead[4519] = 5'h02;
assign _c_doomhead[4520] = 5'h01;
assign _c_doomhead[4521] = 5'h04;
assign _c_doomhead[4522] = 5'h04;
assign _c_doomhead[4523] = 5'h02;
assign _c_doomhead[4524] = 5'h01;
assign _c_doomhead[4525] = 5'h0a;
assign _c_doomhead[4526] = 5'h0f;
assign _c_doomhead[4527] = 5'h14;
assign _c_doomhead[4528] = 5'h19;
assign _c_doomhead[4529] = 5'h1e;
assign _c_doomhead[4530] = 5'h1e;
assign _c_doomhead[4531] = 5'h18;
assign _c_doomhead[4532] = 5'h18;
assign _c_doomhead[4533] = 5'h19;
assign _c_doomhead[4534] = 5'h0d;
assign _c_doomhead[4535] = 5'h0d;
assign _c_doomhead[4536] = 5'h1a;
assign _c_doomhead[4537] = 5'h1c;
assign _c_doomhead[4538] = 5'h0b;
assign _c_doomhead[4539] = 5'h00;
assign _c_doomhead[4540] = 5'h00;
assign _c_doomhead[4541] = 5'h00;
assign _c_doomhead[4542] = 5'h00;
assign _c_doomhead[4543] = 5'h00;
assign _c_doomhead[4544] = 5'h00;
assign _c_doomhead[4545] = 5'h03;
assign _c_doomhead[4546] = 5'h03;
assign _c_doomhead[4547] = 5'h03;
assign _c_doomhead[4548] = 5'h08;
assign _c_doomhead[4549] = 5'h0a;
assign _c_doomhead[4550] = 5'h08;
assign _c_doomhead[4551] = 5'h07;
assign _c_doomhead[4552] = 5'h07;
assign _c_doomhead[4553] = 5'h01;
assign _c_doomhead[4554] = 5'h01;
assign _c_doomhead[4555] = 5'h01;
assign _c_doomhead[4556] = 5'h0b;
assign _c_doomhead[4557] = 5'h0c;
assign _c_doomhead[4558] = 5'h14;
assign _c_doomhead[4559] = 5'h18;
assign _c_doomhead[4560] = 5'h16;
assign _c_doomhead[4561] = 5'h1e;
assign _c_doomhead[4562] = 5'h1e;
assign _c_doomhead[4563] = 5'h16;
assign _c_doomhead[4564] = 5'h16;
assign _c_doomhead[4565] = 5'h16;
assign _c_doomhead[4566] = 5'h16;
assign _c_doomhead[4567] = 5'h16;
assign _c_doomhead[4568] = 5'h1c;
assign _c_doomhead[4569] = 5'h0b;
assign _c_doomhead[4570] = 5'h02;
assign _c_doomhead[4571] = 5'h00;
assign _c_doomhead[4572] = 5'h00;
assign _c_doomhead[4573] = 5'h00;
assign _c_doomhead[4574] = 5'h00;
assign _c_doomhead[4575] = 5'h00;
assign _c_doomhead[4576] = 5'h00;
assign _c_doomhead[4577] = 5'h03;
assign _c_doomhead[4578] = 5'h03;
assign _c_doomhead[4579] = 5'h03;
assign _c_doomhead[4580] = 5'h01;
assign _c_doomhead[4581] = 5'h0a;
assign _c_doomhead[4582] = 5'h0e;
assign _c_doomhead[4583] = 5'h0f;
assign _c_doomhead[4584] = 5'h09;
assign _c_doomhead[4585] = 5'h09;
assign _c_doomhead[4586] = 5'h09;
assign _c_doomhead[4587] = 5'h0b;
assign _c_doomhead[4588] = 5'h0c;
assign _c_doomhead[4589] = 5'h0d;
assign _c_doomhead[4590] = 5'h12;
assign _c_doomhead[4591] = 5'h0f;
assign _c_doomhead[4592] = 5'h09;
assign _c_doomhead[4593] = 5'h03;
assign _c_doomhead[4594] = 5'h03;
assign _c_doomhead[4595] = 5'h07;
assign _c_doomhead[4596] = 5'h0f;
assign _c_doomhead[4597] = 5'h14;
assign _c_doomhead[4598] = 5'h0c;
assign _c_doomhead[4599] = 5'h1e;
assign _c_doomhead[4600] = 5'h02;
assign _c_doomhead[4601] = 5'h10;
assign _c_doomhead[4602] = 5'h10;
assign _c_doomhead[4603] = 5'h00;
assign _c_doomhead[4604] = 5'h00;
assign _c_doomhead[4605] = 5'h00;
assign _c_doomhead[4606] = 5'h00;
assign _c_doomhead[4607] = 5'h00;
assign _c_doomhead[4608] = 5'h00;
assign _c_doomhead[4609] = 5'h03;
assign _c_doomhead[4610] = 5'h03;
assign _c_doomhead[4611] = 5'h03;
assign _c_doomhead[4612] = 5'h04;
assign _c_doomhead[4613] = 5'h07;
assign _c_doomhead[4614] = 5'h0e;
assign _c_doomhead[4615] = 5'h04;
assign _c_doomhead[4616] = 5'h01;
assign _c_doomhead[4617] = 5'h01;
assign _c_doomhead[4618] = 5'h09;
assign _c_doomhead[4619] = 5'h14;
assign _c_doomhead[4620] = 5'h13;
assign _c_doomhead[4621] = 5'h09;
assign _c_doomhead[4622] = 5'h04;
assign _c_doomhead[4623] = 5'h1e;
assign _c_doomhead[4624] = 5'h1c;
assign _c_doomhead[4625] = 5'h17;
assign _c_doomhead[4626] = 5'h03;
assign _c_doomhead[4627] = 5'h1b;
assign _c_doomhead[4628] = 5'h05;
assign _c_doomhead[4629] = 5'h0b;
assign _c_doomhead[4630] = 5'h17;
assign _c_doomhead[4631] = 5'h1a;
assign _c_doomhead[4632] = 5'h17;
assign _c_doomhead[4633] = 5'h10;
assign _c_doomhead[4634] = 5'h00;
assign _c_doomhead[4635] = 5'h00;
assign _c_doomhead[4636] = 5'h00;
assign _c_doomhead[4637] = 5'h00;
assign _c_doomhead[4638] = 5'h00;
assign _c_doomhead[4639] = 5'h00;
assign _c_doomhead[4640] = 5'h00;
assign _c_doomhead[4641] = 5'h00;
assign _c_doomhead[4642] = 5'h03;
assign _c_doomhead[4643] = 5'h03;
assign _c_doomhead[4644] = 5'h03;
assign _c_doomhead[4645] = 5'h04;
assign _c_doomhead[4646] = 5'h0a;
assign _c_doomhead[4647] = 5'h0e;
assign _c_doomhead[4648] = 5'h08;
assign _c_doomhead[4649] = 5'h08;
assign _c_doomhead[4650] = 5'h09;
assign _c_doomhead[4651] = 5'h0c;
assign _c_doomhead[4652] = 5'h0d;
assign _c_doomhead[4653] = 5'h0a;
assign _c_doomhead[4654] = 5'h04;
assign _c_doomhead[4655] = 5'h04;
assign _c_doomhead[4656] = 5'h0c;
assign _c_doomhead[4657] = 5'h1b;
assign _c_doomhead[4658] = 5'h03;
assign _c_doomhead[4659] = 5'h04;
assign _c_doomhead[4660] = 5'h08;
assign _c_doomhead[4661] = 5'h16;
assign _c_doomhead[4662] = 5'h09;
assign _c_doomhead[4663] = 5'h04;
assign _c_doomhead[4664] = 5'h1b;
assign _c_doomhead[4665] = 5'h0b;
assign _c_doomhead[4666] = 5'h00;
assign _c_doomhead[4667] = 5'h00;
assign _c_doomhead[4668] = 5'h00;
assign _c_doomhead[4669] = 5'h00;
assign _c_doomhead[4670] = 5'h00;
assign _c_doomhead[4671] = 5'h00;
assign _c_doomhead[4672] = 5'h00;
assign _c_doomhead[4673] = 5'h00;
assign _c_doomhead[4674] = 5'h03;
assign _c_doomhead[4675] = 5'h03;
assign _c_doomhead[4676] = 5'h03;
assign _c_doomhead[4677] = 5'h0e;
assign _c_doomhead[4678] = 5'h04;
assign _c_doomhead[4679] = 5'h01;
assign _c_doomhead[4680] = 5'h08;
assign _c_doomhead[4681] = 5'h01;
assign _c_doomhead[4682] = 5'h08;
assign _c_doomhead[4683] = 5'h0f;
assign _c_doomhead[4684] = 5'h12;
assign _c_doomhead[4685] = 5'h12;
assign _c_doomhead[4686] = 5'h0d;
assign _c_doomhead[4687] = 5'h07;
assign _c_doomhead[4688] = 5'h02;
assign _c_doomhead[4689] = 5'h02;
assign _c_doomhead[4690] = 5'h02;
assign _c_doomhead[4691] = 5'h08;
assign _c_doomhead[4692] = 5'h07;
assign _c_doomhead[4693] = 5'h14;
assign _c_doomhead[4694] = 5'h0f;
assign _c_doomhead[4695] = 5'h01;
assign _c_doomhead[4696] = 5'h18;
assign _c_doomhead[4697] = 5'h0b;
assign _c_doomhead[4698] = 5'h00;
assign _c_doomhead[4699] = 5'h00;
assign _c_doomhead[4700] = 5'h00;
assign _c_doomhead[4701] = 5'h00;
assign _c_doomhead[4702] = 5'h00;
assign _c_doomhead[4703] = 5'h00;
assign _c_doomhead[4704] = 5'h00;
assign _c_doomhead[4705] = 5'h00;
assign _c_doomhead[4706] = 5'h03;
assign _c_doomhead[4707] = 5'h03;
assign _c_doomhead[4708] = 5'h03;
assign _c_doomhead[4709] = 5'h15;
assign _c_doomhead[4710] = 5'h15;
assign _c_doomhead[4711] = 5'h01;
assign _c_doomhead[4712] = 5'h08;
assign _c_doomhead[4713] = 5'h09;
assign _c_doomhead[4714] = 5'h08;
assign _c_doomhead[4715] = 5'h09;
assign _c_doomhead[4716] = 5'h0c;
assign _c_doomhead[4717] = 5'h18;
assign _c_doomhead[4718] = 5'h16;
assign _c_doomhead[4719] = 5'h16;
assign _c_doomhead[4720] = 5'h0d;
assign _c_doomhead[4721] = 5'h1b;
assign _c_doomhead[4722] = 5'h0d;
assign _c_doomhead[4723] = 5'h01;
assign _c_doomhead[4724] = 5'h07;
assign _c_doomhead[4725] = 5'h14;
assign _c_doomhead[4726] = 5'h0c;
assign _c_doomhead[4727] = 5'h14;
assign _c_doomhead[4728] = 5'h18;
assign _c_doomhead[4729] = 5'h07;
assign _c_doomhead[4730] = 5'h00;
assign _c_doomhead[4731] = 5'h00;
assign _c_doomhead[4732] = 5'h00;
assign _c_doomhead[4733] = 5'h00;
assign _c_doomhead[4734] = 5'h00;
assign _c_doomhead[4735] = 5'h00;
assign _c_doomhead[4736] = 5'h00;
assign _c_doomhead[4737] = 5'h00;
assign _c_doomhead[4738] = 5'h03;
assign _c_doomhead[4739] = 5'h03;
assign _c_doomhead[4740] = 5'h03;
assign _c_doomhead[4741] = 5'h15;
assign _c_doomhead[4742] = 5'h15;
assign _c_doomhead[4743] = 5'h08;
assign _c_doomhead[4744] = 5'h01;
assign _c_doomhead[4745] = 5'h0f;
assign _c_doomhead[4746] = 5'h08;
assign _c_doomhead[4747] = 5'h08;
assign _c_doomhead[4748] = 5'h0a;
assign _c_doomhead[4749] = 5'h18;
assign _c_doomhead[4750] = 5'h16;
assign _c_doomhead[4751] = 5'h14;
assign _c_doomhead[4752] = 5'h1b;
assign _c_doomhead[4753] = 5'h1b;
assign _c_doomhead[4754] = 5'h0b;
assign _c_doomhead[4755] = 5'h12;
assign _c_doomhead[4756] = 5'h0f;
assign _c_doomhead[4757] = 5'h18;
assign _c_doomhead[4758] = 5'h14;
assign _c_doomhead[4759] = 5'h14;
assign _c_doomhead[4760] = 5'h0d;
assign _c_doomhead[4761] = 5'h08;
assign _c_doomhead[4762] = 5'h00;
assign _c_doomhead[4763] = 5'h00;
assign _c_doomhead[4764] = 5'h00;
assign _c_doomhead[4765] = 5'h00;
assign _c_doomhead[4766] = 5'h00;
assign _c_doomhead[4767] = 5'h00;
assign _c_doomhead[4768] = 5'h00;
assign _c_doomhead[4769] = 5'h00;
assign _c_doomhead[4770] = 5'h00;
assign _c_doomhead[4771] = 5'h03;
assign _c_doomhead[4772] = 5'h03;
assign _c_doomhead[4773] = 5'h01;
assign _c_doomhead[4774] = 5'h15;
assign _c_doomhead[4775] = 5'h07;
assign _c_doomhead[4776] = 5'h09;
assign _c_doomhead[4777] = 5'h0f;
assign _c_doomhead[4778] = 5'h08;
assign _c_doomhead[4779] = 5'h08;
assign _c_doomhead[4780] = 5'h0f;
assign _c_doomhead[4781] = 5'h19;
assign _c_doomhead[4782] = 5'h16;
assign _c_doomhead[4783] = 5'h1e;
assign _c_doomhead[4784] = 5'h1c;
assign _c_doomhead[4785] = 5'h08;
assign _c_doomhead[4786] = 5'h1c;
assign _c_doomhead[4787] = 5'h06;
assign _c_doomhead[4788] = 5'h0a;
assign _c_doomhead[4789] = 5'h18;
assign _c_doomhead[4790] = 5'h0f;
assign _c_doomhead[4791] = 5'h0d;
assign _c_doomhead[4792] = 5'h01;
assign _c_doomhead[4793] = 5'h00;
assign _c_doomhead[4794] = 5'h00;
assign _c_doomhead[4795] = 5'h00;
assign _c_doomhead[4796] = 5'h00;
assign _c_doomhead[4797] = 5'h00;
assign _c_doomhead[4798] = 5'h00;
assign _c_doomhead[4799] = 5'h00;
assign _c_doomhead[4800] = 5'h00;
assign _c_doomhead[4801] = 5'h00;
assign _c_doomhead[4802] = 5'h00;
assign _c_doomhead[4803] = 5'h00;
assign _c_doomhead[4804] = 5'h15;
assign _c_doomhead[4805] = 5'h01;
assign _c_doomhead[4806] = 5'h01;
assign _c_doomhead[4807] = 5'h07;
assign _c_doomhead[4808] = 5'h07;
assign _c_doomhead[4809] = 5'h0b;
assign _c_doomhead[4810] = 5'h01;
assign _c_doomhead[4811] = 5'h08;
assign _c_doomhead[4812] = 5'h0c;
assign _c_doomhead[4813] = 5'h19;
assign _c_doomhead[4814] = 5'h0c;
assign _c_doomhead[4815] = 5'h1c;
assign _c_doomhead[4816] = 5'h0c;
assign _c_doomhead[4817] = 5'h09;
assign _c_doomhead[4818] = 5'h1c;
assign _c_doomhead[4819] = 5'h1c;
assign _c_doomhead[4820] = 5'h04;
assign _c_doomhead[4821] = 5'h0a;
assign _c_doomhead[4822] = 5'h01;
assign _c_doomhead[4823] = 5'h0b;
assign _c_doomhead[4824] = 5'h04;
assign _c_doomhead[4825] = 5'h00;
assign _c_doomhead[4826] = 5'h00;
assign _c_doomhead[4827] = 5'h00;
assign _c_doomhead[4828] = 5'h00;
assign _c_doomhead[4829] = 5'h00;
assign _c_doomhead[4830] = 5'h00;
assign _c_doomhead[4831] = 5'h00;
assign _c_doomhead[4832] = 5'h00;
assign _c_doomhead[4833] = 5'h00;
assign _c_doomhead[4834] = 5'h00;
assign _c_doomhead[4835] = 5'h00;
assign _c_doomhead[4836] = 5'h00;
assign _c_doomhead[4837] = 5'h07;
assign _c_doomhead[4838] = 5'h01;
assign _c_doomhead[4839] = 5'h15;
assign _c_doomhead[4840] = 5'h07;
assign _c_doomhead[4841] = 5'h07;
assign _c_doomhead[4842] = 5'h07;
assign _c_doomhead[4843] = 5'h01;
assign _c_doomhead[4844] = 5'h0c;
assign _c_doomhead[4845] = 5'h12;
assign _c_doomhead[4846] = 5'h09;
assign _c_doomhead[4847] = 5'h1c;
assign _c_doomhead[4848] = 5'h14;
assign _c_doomhead[4849] = 5'h0c;
assign _c_doomhead[4850] = 5'h1c;
assign _c_doomhead[4851] = 5'h1c;
assign _c_doomhead[4852] = 5'h03;
assign _c_doomhead[4853] = 5'h1a;
assign _c_doomhead[4854] = 5'h1a;
assign _c_doomhead[4855] = 5'h07;
assign _c_doomhead[4856] = 5'h00;
assign _c_doomhead[4857] = 5'h00;
assign _c_doomhead[4858] = 5'h00;
assign _c_doomhead[4859] = 5'h00;
assign _c_doomhead[4860] = 5'h00;
assign _c_doomhead[4861] = 5'h00;
assign _c_doomhead[4862] = 5'h00;
assign _c_doomhead[4863] = 5'h00;
assign _c_doomhead[4864] = 5'h00;
assign _c_doomhead[4865] = 5'h00;
assign _c_doomhead[4866] = 5'h00;
assign _c_doomhead[4867] = 5'h00;
assign _c_doomhead[4868] = 5'h00;
assign _c_doomhead[4869] = 5'h00;
assign _c_doomhead[4870] = 5'h01;
assign _c_doomhead[4871] = 5'h02;
assign _c_doomhead[4872] = 5'h08;
assign _c_doomhead[4873] = 5'h07;
assign _c_doomhead[4874] = 5'h07;
assign _c_doomhead[4875] = 5'h01;
assign _c_doomhead[4876] = 5'h0f;
assign _c_doomhead[4877] = 5'h14;
assign _c_doomhead[4878] = 5'h09;
assign _c_doomhead[4879] = 5'h1c;
assign _c_doomhead[4880] = 5'h0c;
assign _c_doomhead[4881] = 5'h19;
assign _c_doomhead[4882] = 5'h1e;
assign _c_doomhead[4883] = 5'h1e;
assign _c_doomhead[4884] = 5'h1d;
assign _c_doomhead[4885] = 5'h1d;
assign _c_doomhead[4886] = 5'h1b;
assign _c_doomhead[4887] = 5'h01;
assign _c_doomhead[4888] = 5'h00;
assign _c_doomhead[4889] = 5'h00;
assign _c_doomhead[4890] = 5'h00;
assign _c_doomhead[4891] = 5'h00;
assign _c_doomhead[4892] = 5'h00;
assign _c_doomhead[4893] = 5'h00;
assign _c_doomhead[4894] = 5'h00;
assign _c_doomhead[4895] = 5'h00;
assign _c_doomhead[4896] = 5'h00;
assign _c_doomhead[4897] = 5'h00;
assign _c_doomhead[4898] = 5'h00;
assign _c_doomhead[4899] = 5'h00;
assign _c_doomhead[4900] = 5'h00;
assign _c_doomhead[4901] = 5'h00;
assign _c_doomhead[4902] = 5'h00;
assign _c_doomhead[4903] = 5'h04;
assign _c_doomhead[4904] = 5'h02;
assign _c_doomhead[4905] = 5'h15;
assign _c_doomhead[4906] = 5'h07;
assign _c_doomhead[4907] = 5'h0b;
assign _c_doomhead[4908] = 5'h0f;
assign _c_doomhead[4909] = 5'h0c;
assign _c_doomhead[4910] = 5'h0f;
assign _c_doomhead[4911] = 5'h1b;
assign _c_doomhead[4912] = 5'h09;
assign _c_doomhead[4913] = 5'h1d;
assign _c_doomhead[4914] = 5'h1b;
assign _c_doomhead[4915] = 5'h1c;
assign _c_doomhead[4916] = 5'h1c;
assign _c_doomhead[4917] = 5'h1c;
assign _c_doomhead[4918] = 5'h09;
assign _c_doomhead[4919] = 5'h04;
assign _c_doomhead[4920] = 5'h00;
assign _c_doomhead[4921] = 5'h00;
assign _c_doomhead[4922] = 5'h00;
assign _c_doomhead[4923] = 5'h00;
assign _c_doomhead[4924] = 5'h00;
assign _c_doomhead[4925] = 5'h00;
assign _c_doomhead[4926] = 5'h00;
assign _c_doomhead[4927] = 5'h00;
assign _c_doomhead[4928] = 5'h00;
assign _c_doomhead[4929] = 5'h00;
assign _c_doomhead[4930] = 5'h00;
assign _c_doomhead[4931] = 5'h00;
assign _c_doomhead[4932] = 5'h00;
assign _c_doomhead[4933] = 5'h00;
assign _c_doomhead[4934] = 5'h00;
assign _c_doomhead[4935] = 5'h00;
assign _c_doomhead[4936] = 5'h04;
assign _c_doomhead[4937] = 5'h15;
assign _c_doomhead[4938] = 5'h07;
assign _c_doomhead[4939] = 5'h0f;
assign _c_doomhead[4940] = 5'h0f;
assign _c_doomhead[4941] = 5'h13;
assign _c_doomhead[4942] = 5'h1e;
assign _c_doomhead[4943] = 5'h1e;
assign _c_doomhead[4944] = 5'h0b;
assign _c_doomhead[4945] = 5'h0c;
assign _c_doomhead[4946] = 5'h1e;
assign _c_doomhead[4947] = 5'h1e;
assign _c_doomhead[4948] = 5'h0c;
assign _c_doomhead[4949] = 5'h0f;
assign _c_doomhead[4950] = 5'h1d;
assign _c_doomhead[4951] = 5'h00;
assign _c_doomhead[4952] = 5'h00;
assign _c_doomhead[4953] = 5'h00;
assign _c_doomhead[4954] = 5'h00;
assign _c_doomhead[4955] = 5'h00;
assign _c_doomhead[4956] = 5'h00;
assign _c_doomhead[4957] = 5'h00;
assign _c_doomhead[4958] = 5'h00;
assign _c_doomhead[4959] = 5'h00;
assign _c_doomhead[4960] = 5'h00;
assign _c_doomhead[4961] = 5'h00;
assign _c_doomhead[4962] = 5'h00;
assign _c_doomhead[4963] = 5'h00;
assign _c_doomhead[4964] = 5'h00;
assign _c_doomhead[4965] = 5'h00;
assign _c_doomhead[4966] = 5'h00;
assign _c_doomhead[4967] = 5'h00;
assign _c_doomhead[4968] = 5'h00;
assign _c_doomhead[4969] = 5'h05;
assign _c_doomhead[4970] = 5'h02;
assign _c_doomhead[4971] = 5'h07;
assign _c_doomhead[4972] = 5'h0b;
assign _c_doomhead[4973] = 5'h0f;
assign _c_doomhead[4974] = 5'h1b;
assign _c_doomhead[4975] = 5'h0b;
assign _c_doomhead[4976] = 5'h07;
assign _c_doomhead[4977] = 5'h07;
assign _c_doomhead[4978] = 5'h1c;
assign _c_doomhead[4979] = 5'h1c;
assign _c_doomhead[4980] = 5'h1c;
assign _c_doomhead[4981] = 5'h1a;
assign _c_doomhead[4982] = 5'h01;
assign _c_doomhead[4983] = 5'h00;
assign _c_doomhead[4984] = 5'h00;
assign _c_doomhead[4985] = 5'h00;
assign _c_doomhead[4986] = 5'h00;
assign _c_doomhead[4987] = 5'h00;
assign _c_doomhead[4988] = 5'h00;
assign _c_doomhead[4989] = 5'h00;
assign _c_doomhead[4990] = 5'h00;
assign _c_doomhead[4991] = 5'h00;
assign _c_doomhead[4992] = 5'h00;
assign _c_doomhead[4993] = 5'h00;
assign _c_doomhead[4994] = 5'h00;
assign _c_doomhead[4995] = 5'h00;
assign _c_doomhead[4996] = 5'h00;
assign _c_doomhead[4997] = 5'h00;
assign _c_doomhead[4998] = 5'h00;
assign _c_doomhead[4999] = 5'h00;
assign _c_doomhead[5000] = 5'h00;
assign _c_doomhead[5001] = 5'h00;
assign _c_doomhead[5002] = 5'h00;
assign _c_doomhead[5003] = 5'h05;
assign _c_doomhead[5004] = 5'h15;
assign _c_doomhead[5005] = 5'h07;
assign _c_doomhead[5006] = 5'h1b;
assign _c_doomhead[5007] = 5'h0f;
assign _c_doomhead[5008] = 5'h0f;
assign _c_doomhead[5009] = 5'h0c;
assign _c_doomhead[5010] = 5'h1b;
assign _c_doomhead[5011] = 5'h1b;
assign _c_doomhead[5012] = 5'h1a;
assign _c_doomhead[5013] = 5'h01;
assign _c_doomhead[5014] = 5'h04;
assign _c_doomhead[5015] = 5'h00;
assign _c_doomhead[5016] = 5'h00;
assign _c_doomhead[5017] = 5'h00;
assign _c_doomhead[5018] = 5'h00;
assign _c_doomhead[5019] = 5'h00;
assign _c_doomhead[5020] = 5'h00;
assign _c_doomhead[5021] = 5'h00;
assign _c_doomhead[5022] = 5'h00;
assign _c_doomhead[5023] = 5'h00;
assign _c_doomhead[5024] = 5'h00;
assign _c_doomhead[5025] = 5'h00;
assign _c_doomhead[5026] = 5'h00;
assign _c_doomhead[5027] = 5'h00;
assign _c_doomhead[5028] = 5'h00;
assign _c_doomhead[5029] = 5'h00;
assign _c_doomhead[5030] = 5'h00;
assign _c_doomhead[5031] = 5'h00;
assign _c_doomhead[5032] = 5'h00;
assign _c_doomhead[5033] = 5'h00;
assign _c_doomhead[5034] = 5'h00;
assign _c_doomhead[5035] = 5'h00;
assign _c_doomhead[5036] = 5'h05;
assign _c_doomhead[5037] = 5'h05;
assign _c_doomhead[5038] = 5'h1a;
assign _c_doomhead[5039] = 5'h01;
assign _c_doomhead[5040] = 5'h09;
assign _c_doomhead[5041] = 5'h1d;
assign _c_doomhead[5042] = 5'h1c;
assign _c_doomhead[5043] = 5'h1c;
assign _c_doomhead[5044] = 5'h1a;
assign _c_doomhead[5045] = 5'h04;
assign _c_doomhead[5046] = 5'h00;
assign _c_doomhead[5047] = 5'h00;
assign _c_doomhead[5048] = 5'h00;
assign _c_doomhead[5049] = 5'h00;
assign _c_doomhead[5050] = 5'h00;
assign _c_doomhead[5051] = 5'h00;
assign _c_doomhead[5052] = 5'h00;
assign _c_doomhead[5053] = 5'h00;
assign _c_doomhead[5054] = 5'h00;
assign _c_doomhead[5055] = 5'h00;
assign _c_doomhead[5056] = 5'h00;
assign _c_doomhead[5057] = 5'h00;
assign _c_doomhead[5058] = 5'h00;
assign _c_doomhead[5059] = 5'h00;
assign _c_doomhead[5060] = 5'h00;
assign _c_doomhead[5061] = 5'h00;
assign _c_doomhead[5062] = 5'h00;
assign _c_doomhead[5063] = 5'h00;
assign _c_doomhead[5064] = 5'h00;
assign _c_doomhead[5065] = 5'h00;
assign _c_doomhead[5066] = 5'h00;
assign _c_doomhead[5067] = 5'h00;
assign _c_doomhead[5068] = 5'h00;
assign _c_doomhead[5069] = 5'h00;
assign _c_doomhead[5070] = 5'h00;
assign _c_doomhead[5071] = 5'h00;
assign _c_doomhead[5072] = 5'h00;
assign _c_doomhead[5073] = 5'h00;
assign _c_doomhead[5074] = 5'h00;
assign _c_doomhead[5075] = 5'h00;
assign _c_doomhead[5076] = 5'h00;
assign _c_doomhead[5077] = 5'h00;
assign _c_doomhead[5078] = 5'h00;
assign _c_doomhead[5079] = 5'h00;
assign _c_doomhead[5080] = 5'h00;
assign _c_doomhead[5081] = 5'h00;
assign _c_doomhead[5082] = 5'h00;
assign _c_doomhead[5083] = 5'h00;
assign _c_doomhead[5084] = 5'h00;
assign _c_doomhead[5085] = 5'h00;
assign _c_doomhead[5086] = 5'h00;
assign _c_doomhead[5087] = 5'h00;
assign _c_doomhead[5088] = 5'h00;
assign _c_doomhead[5089] = 5'h00;
assign _c_doomhead[5090] = 5'h00;
assign _c_doomhead[5091] = 5'h00;
assign _c_doomhead[5092] = 5'h00;
assign _c_doomhead[5093] = 5'h00;
assign _c_doomhead[5094] = 5'h00;
assign _c_doomhead[5095] = 5'h00;
assign _c_doomhead[5096] = 5'h00;
assign _c_doomhead[5097] = 5'h00;
assign _c_doomhead[5098] = 5'h00;
assign _c_doomhead[5099] = 5'h00;
assign _c_doomhead[5100] = 5'h00;
assign _c_doomhead[5101] = 5'h00;
assign _c_doomhead[5102] = 5'h00;
assign _c_doomhead[5103] = 5'h00;
assign _c_doomhead[5104] = 5'h00;
assign _c_doomhead[5105] = 5'h00;
assign _c_doomhead[5106] = 5'h00;
assign _c_doomhead[5107] = 5'h00;
assign _c_doomhead[5108] = 5'h00;
assign _c_doomhead[5109] = 5'h00;
assign _c_doomhead[5110] = 5'h00;
assign _c_doomhead[5111] = 5'h00;
assign _c_doomhead[5112] = 5'h00;
assign _c_doomhead[5113] = 5'h00;
assign _c_doomhead[5114] = 5'h00;
assign _c_doomhead[5115] = 5'h00;
assign _c_doomhead[5116] = 5'h00;
assign _c_doomhead[5117] = 5'h00;
assign _c_doomhead[5118] = 5'h00;
assign _c_doomhead[5119] = 5'h00;
assign _c_doomhead[5120] = 5'h00;
assign _c_doomhead[5121] = 5'h00;
assign _c_doomhead[5122] = 5'h00;
assign _c_doomhead[5123] = 5'h00;
assign _c_doomhead[5124] = 5'h00;
assign _c_doomhead[5125] = 5'h00;
assign _c_doomhead[5126] = 5'h00;
assign _c_doomhead[5127] = 5'h00;
assign _c_doomhead[5128] = 5'h05;
assign _c_doomhead[5129] = 5'h02;
assign _c_doomhead[5130] = 5'h02;
assign _c_doomhead[5131] = 5'h04;
assign _c_doomhead[5132] = 5'h06;
assign _c_doomhead[5133] = 5'h06;
assign _c_doomhead[5134] = 5'h06;
assign _c_doomhead[5135] = 5'h06;
assign _c_doomhead[5136] = 5'h06;
assign _c_doomhead[5137] = 5'h06;
assign _c_doomhead[5138] = 5'h04;
assign _c_doomhead[5139] = 5'h02;
assign _c_doomhead[5140] = 5'h02;
assign _c_doomhead[5141] = 5'h05;
assign _c_doomhead[5142] = 5'h00;
assign _c_doomhead[5143] = 5'h00;
assign _c_doomhead[5144] = 5'h00;
assign _c_doomhead[5145] = 5'h00;
assign _c_doomhead[5146] = 5'h00;
assign _c_doomhead[5147] = 5'h00;
assign _c_doomhead[5148] = 5'h00;
assign _c_doomhead[5149] = 5'h00;
assign _c_doomhead[5150] = 5'h00;
assign _c_doomhead[5151] = 5'h00;
assign _c_doomhead[5152] = 5'h00;
assign _c_doomhead[5153] = 5'h00;
assign _c_doomhead[5154] = 5'h00;
assign _c_doomhead[5155] = 5'h00;
assign _c_doomhead[5156] = 5'h00;
assign _c_doomhead[5157] = 5'h00;
assign _c_doomhead[5158] = 5'h03;
assign _c_doomhead[5159] = 5'h02;
assign _c_doomhead[5160] = 5'h0e;
assign _c_doomhead[5161] = 5'h02;
assign _c_doomhead[5162] = 5'h04;
assign _c_doomhead[5163] = 5'h06;
assign _c_doomhead[5164] = 5'h01;
assign _c_doomhead[5165] = 5'h07;
assign _c_doomhead[5166] = 5'h07;
assign _c_doomhead[5167] = 5'h07;
assign _c_doomhead[5168] = 5'h07;
assign _c_doomhead[5169] = 5'h01;
assign _c_doomhead[5170] = 5'h06;
assign _c_doomhead[5171] = 5'h04;
assign _c_doomhead[5172] = 5'h02;
assign _c_doomhead[5173] = 5'h0e;
assign _c_doomhead[5174] = 5'h02;
assign _c_doomhead[5175] = 5'h03;
assign _c_doomhead[5176] = 5'h00;
assign _c_doomhead[5177] = 5'h00;
assign _c_doomhead[5178] = 5'h00;
assign _c_doomhead[5179] = 5'h00;
assign _c_doomhead[5180] = 5'h00;
assign _c_doomhead[5181] = 5'h00;
assign _c_doomhead[5182] = 5'h00;
assign _c_doomhead[5183] = 5'h00;
assign _c_doomhead[5184] = 5'h00;
assign _c_doomhead[5185] = 5'h00;
assign _c_doomhead[5186] = 5'h00;
assign _c_doomhead[5187] = 5'h00;
assign _c_doomhead[5188] = 5'h00;
assign _c_doomhead[5189] = 5'h03;
assign _c_doomhead[5190] = 5'h0e;
assign _c_doomhead[5191] = 5'h04;
assign _c_doomhead[5192] = 5'h01;
assign _c_doomhead[5193] = 5'h01;
assign _c_doomhead[5194] = 5'h09;
assign _c_doomhead[5195] = 5'h09;
assign _c_doomhead[5196] = 5'h0b;
assign _c_doomhead[5197] = 5'h0b;
assign _c_doomhead[5198] = 5'h0f;
assign _c_doomhead[5199] = 5'h0a;
assign _c_doomhead[5200] = 5'h0b;
assign _c_doomhead[5201] = 5'h07;
assign _c_doomhead[5202] = 5'h01;
assign _c_doomhead[5203] = 5'h08;
assign _c_doomhead[5204] = 5'h06;
assign _c_doomhead[5205] = 5'h06;
assign _c_doomhead[5206] = 5'h04;
assign _c_doomhead[5207] = 5'h05;
assign _c_doomhead[5208] = 5'h03;
assign _c_doomhead[5209] = 5'h00;
assign _c_doomhead[5210] = 5'h00;
assign _c_doomhead[5211] = 5'h00;
assign _c_doomhead[5212] = 5'h00;
assign _c_doomhead[5213] = 5'h00;
assign _c_doomhead[5214] = 5'h00;
assign _c_doomhead[5215] = 5'h00;
assign _c_doomhead[5216] = 5'h00;
assign _c_doomhead[5217] = 5'h00;
assign _c_doomhead[5218] = 5'h00;
assign _c_doomhead[5219] = 5'h00;
assign _c_doomhead[5220] = 5'h00;
assign _c_doomhead[5221] = 5'h03;
assign _c_doomhead[5222] = 5'h05;
assign _c_doomhead[5223] = 5'h01;
assign _c_doomhead[5224] = 5'h01;
assign _c_doomhead[5225] = 5'h09;
assign _c_doomhead[5226] = 5'h09;
assign _c_doomhead[5227] = 5'h0a;
assign _c_doomhead[5228] = 5'h0a;
assign _c_doomhead[5229] = 5'h0f;
assign _c_doomhead[5230] = 5'h0f;
assign _c_doomhead[5231] = 5'h0f;
assign _c_doomhead[5232] = 5'h0f;
assign _c_doomhead[5233] = 5'h0a;
assign _c_doomhead[5234] = 5'h09;
assign _c_doomhead[5235] = 5'h01;
assign _c_doomhead[5236] = 5'h01;
assign _c_doomhead[5237] = 5'h08;
assign _c_doomhead[5238] = 5'h04;
assign _c_doomhead[5239] = 5'h05;
assign _c_doomhead[5240] = 5'h11;
assign _c_doomhead[5241] = 5'h00;
assign _c_doomhead[5242] = 5'h00;
assign _c_doomhead[5243] = 5'h00;
assign _c_doomhead[5244] = 5'h00;
assign _c_doomhead[5245] = 5'h00;
assign _c_doomhead[5246] = 5'h00;
assign _c_doomhead[5247] = 5'h00;
assign _c_doomhead[5248] = 5'h00;
assign _c_doomhead[5249] = 5'h00;
assign _c_doomhead[5250] = 5'h00;
assign _c_doomhead[5251] = 5'h00;
assign _c_doomhead[5252] = 5'h11;
assign _c_doomhead[5253] = 5'h03;
assign _c_doomhead[5254] = 5'h0e;
assign _c_doomhead[5255] = 5'h02;
assign _c_doomhead[5256] = 5'h06;
assign _c_doomhead[5257] = 5'h01;
assign _c_doomhead[5258] = 5'h07;
assign _c_doomhead[5259] = 5'h0f;
assign _c_doomhead[5260] = 5'h13;
assign _c_doomhead[5261] = 5'h0c;
assign _c_doomhead[5262] = 5'h09;
assign _c_doomhead[5263] = 5'h0a;
assign _c_doomhead[5264] = 5'h07;
assign _c_doomhead[5265] = 5'h07;
assign _c_doomhead[5266] = 5'h07;
assign _c_doomhead[5267] = 5'h01;
assign _c_doomhead[5268] = 5'h01;
assign _c_doomhead[5269] = 5'h06;
assign _c_doomhead[5270] = 5'h06;
assign _c_doomhead[5271] = 5'h0e;
assign _c_doomhead[5272] = 5'h11;
assign _c_doomhead[5273] = 5'h11;
assign _c_doomhead[5274] = 5'h00;
assign _c_doomhead[5275] = 5'h00;
assign _c_doomhead[5276] = 5'h00;
assign _c_doomhead[5277] = 5'h00;
assign _c_doomhead[5278] = 5'h00;
assign _c_doomhead[5279] = 5'h00;
assign _c_doomhead[5280] = 5'h00;
assign _c_doomhead[5281] = 5'h00;
assign _c_doomhead[5282] = 5'h00;
assign _c_doomhead[5283] = 5'h00;
assign _c_doomhead[5284] = 5'h11;
assign _c_doomhead[5285] = 5'h11;
assign _c_doomhead[5286] = 5'h03;
assign _c_doomhead[5287] = 5'h06;
assign _c_doomhead[5288] = 5'h08;
assign _c_doomhead[5289] = 5'h06;
assign _c_doomhead[5290] = 5'h01;
assign _c_doomhead[5291] = 5'h07;
assign _c_doomhead[5292] = 5'h0a;
assign _c_doomhead[5293] = 5'h0a;
assign _c_doomhead[5294] = 5'h0b;
assign _c_doomhead[5295] = 5'h01;
assign _c_doomhead[5296] = 5'h09;
assign _c_doomhead[5297] = 5'h09;
assign _c_doomhead[5298] = 5'h06;
assign _c_doomhead[5299] = 5'h06;
assign _c_doomhead[5300] = 5'h06;
assign _c_doomhead[5301] = 5'h02;
assign _c_doomhead[5302] = 5'h0e;
assign _c_doomhead[5303] = 5'h03;
assign _c_doomhead[5304] = 5'h03;
assign _c_doomhead[5305] = 5'h11;
assign _c_doomhead[5306] = 5'h00;
assign _c_doomhead[5307] = 5'h00;
assign _c_doomhead[5308] = 5'h00;
assign _c_doomhead[5309] = 5'h00;
assign _c_doomhead[5310] = 5'h00;
assign _c_doomhead[5311] = 5'h00;
assign _c_doomhead[5312] = 5'h00;
assign _c_doomhead[5313] = 5'h00;
assign _c_doomhead[5314] = 5'h00;
assign _c_doomhead[5315] = 5'h00;
assign _c_doomhead[5316] = 5'h11;
assign _c_doomhead[5317] = 5'h11;
assign _c_doomhead[5318] = 5'h11;
assign _c_doomhead[5319] = 5'h02;
assign _c_doomhead[5320] = 5'h06;
assign _c_doomhead[5321] = 5'h02;
assign _c_doomhead[5322] = 5'h0e;
assign _c_doomhead[5323] = 5'h06;
assign _c_doomhead[5324] = 5'h0a;
assign _c_doomhead[5325] = 5'h01;
assign _c_doomhead[5326] = 5'h06;
assign _c_doomhead[5327] = 5'h04;
assign _c_doomhead[5328] = 5'h0a;
assign _c_doomhead[5329] = 5'h01;
assign _c_doomhead[5330] = 5'h02;
assign _c_doomhead[5331] = 5'h03;
assign _c_doomhead[5332] = 5'h02;
assign _c_doomhead[5333] = 5'h05;
assign _c_doomhead[5334] = 5'h03;
assign _c_doomhead[5335] = 5'h11;
assign _c_doomhead[5336] = 5'h03;
assign _c_doomhead[5337] = 5'h11;
assign _c_doomhead[5338] = 5'h00;
assign _c_doomhead[5339] = 5'h00;
assign _c_doomhead[5340] = 5'h00;
assign _c_doomhead[5341] = 5'h00;
assign _c_doomhead[5342] = 5'h00;
assign _c_doomhead[5343] = 5'h00;
assign _c_doomhead[5344] = 5'h00;
assign _c_doomhead[5345] = 5'h00;
assign _c_doomhead[5346] = 5'h00;
assign _c_doomhead[5347] = 5'h00;
assign _c_doomhead[5348] = 5'h11;
assign _c_doomhead[5349] = 5'h03;
assign _c_doomhead[5350] = 5'h03;
assign _c_doomhead[5351] = 5'h05;
assign _c_doomhead[5352] = 5'h0e;
assign _c_doomhead[5353] = 5'h02;
assign _c_doomhead[5354] = 5'h0e;
assign _c_doomhead[5355] = 5'h06;
assign _c_doomhead[5356] = 5'h01;
assign _c_doomhead[5357] = 5'h01;
assign _c_doomhead[5358] = 5'h06;
assign _c_doomhead[5359] = 5'h04;
assign _c_doomhead[5360] = 5'h01;
assign _c_doomhead[5361] = 5'h06;
assign _c_doomhead[5362] = 5'h02;
assign _c_doomhead[5363] = 5'h03;
assign _c_doomhead[5364] = 5'h10;
assign _c_doomhead[5365] = 5'h02;
assign _c_doomhead[5366] = 5'h11;
assign _c_doomhead[5367] = 5'h03;
assign _c_doomhead[5368] = 5'h03;
assign _c_doomhead[5369] = 5'h11;
assign _c_doomhead[5370] = 5'h00;
assign _c_doomhead[5371] = 5'h00;
assign _c_doomhead[5372] = 5'h00;
assign _c_doomhead[5373] = 5'h00;
assign _c_doomhead[5374] = 5'h00;
assign _c_doomhead[5375] = 5'h00;
assign _c_doomhead[5376] = 5'h00;
assign _c_doomhead[5377] = 5'h00;
assign _c_doomhead[5378] = 5'h00;
assign _c_doomhead[5379] = 5'h00;
assign _c_doomhead[5380] = 5'h11;
assign _c_doomhead[5381] = 5'h03;
assign _c_doomhead[5382] = 5'h11;
assign _c_doomhead[5383] = 5'h05;
assign _c_doomhead[5384] = 5'h1c;
assign _c_doomhead[5385] = 5'h1c;
assign _c_doomhead[5386] = 5'h05;
assign _c_doomhead[5387] = 5'h04;
assign _c_doomhead[5388] = 5'h01;
assign _c_doomhead[5389] = 5'h08;
assign _c_doomhead[5390] = 5'h03;
assign _c_doomhead[5391] = 5'h02;
assign _c_doomhead[5392] = 5'h06;
assign _c_doomhead[5393] = 5'h06;
assign _c_doomhead[5394] = 5'h05;
assign _c_doomhead[5395] = 5'h03;
assign _c_doomhead[5396] = 5'h05;
assign _c_doomhead[5397] = 5'h04;
assign _c_doomhead[5398] = 5'h0e;
assign _c_doomhead[5399] = 5'h05;
assign _c_doomhead[5400] = 5'h05;
assign _c_doomhead[5401] = 5'h11;
assign _c_doomhead[5402] = 5'h00;
assign _c_doomhead[5403] = 5'h00;
assign _c_doomhead[5404] = 5'h00;
assign _c_doomhead[5405] = 5'h00;
assign _c_doomhead[5406] = 5'h00;
assign _c_doomhead[5407] = 5'h00;
assign _c_doomhead[5408] = 5'h00;
assign _c_doomhead[5409] = 5'h00;
assign _c_doomhead[5410] = 5'h00;
assign _c_doomhead[5411] = 5'h00;
assign _c_doomhead[5412] = 5'h11;
assign _c_doomhead[5413] = 5'h03;
assign _c_doomhead[5414] = 5'h02;
assign _c_doomhead[5415] = 5'h1c;
assign _c_doomhead[5416] = 5'h1b;
assign _c_doomhead[5417] = 5'h1c;
assign _c_doomhead[5418] = 5'h05;
assign _c_doomhead[5419] = 5'h02;
assign _c_doomhead[5420] = 5'h08;
assign _c_doomhead[5421] = 5'h03;
assign _c_doomhead[5422] = 5'h07;
assign _c_doomhead[5423] = 5'h02;
assign _c_doomhead[5424] = 5'h06;
assign _c_doomhead[5425] = 5'h02;
assign _c_doomhead[5426] = 5'h03;
assign _c_doomhead[5427] = 5'h1b;
assign _c_doomhead[5428] = 5'h1c;
assign _c_doomhead[5429] = 5'h04;
assign _c_doomhead[5430] = 5'h01;
assign _c_doomhead[5431] = 5'h0e;
assign _c_doomhead[5432] = 5'h05;
assign _c_doomhead[5433] = 5'h11;
assign _c_doomhead[5434] = 5'h00;
assign _c_doomhead[5435] = 5'h00;
assign _c_doomhead[5436] = 5'h00;
assign _c_doomhead[5437] = 5'h00;
assign _c_doomhead[5438] = 5'h00;
assign _c_doomhead[5439] = 5'h00;
assign _c_doomhead[5440] = 5'h00;
assign _c_doomhead[5441] = 5'h00;
assign _c_doomhead[5442] = 5'h00;
assign _c_doomhead[5443] = 5'h00;
assign _c_doomhead[5444] = 5'h11;
assign _c_doomhead[5445] = 5'h05;
assign _c_doomhead[5446] = 5'h02;
assign _c_doomhead[5447] = 5'h02;
assign _c_doomhead[5448] = 5'h1c;
assign _c_doomhead[5449] = 5'h1c;
assign _c_doomhead[5450] = 5'h0a;
assign _c_doomhead[5451] = 5'h03;
assign _c_doomhead[5452] = 5'h0e;
assign _c_doomhead[5453] = 5'h03;
assign _c_doomhead[5454] = 5'h09;
assign _c_doomhead[5455] = 5'h03;
assign _c_doomhead[5456] = 5'h06;
assign _c_doomhead[5457] = 5'h03;
assign _c_doomhead[5458] = 5'h04;
assign _c_doomhead[5459] = 5'h1c;
assign _c_doomhead[5460] = 5'h1c;
assign _c_doomhead[5461] = 5'h08;
assign _c_doomhead[5462] = 5'h0b;
assign _c_doomhead[5463] = 5'h01;
assign _c_doomhead[5464] = 5'h05;
assign _c_doomhead[5465] = 5'h11;
assign _c_doomhead[5466] = 5'h00;
assign _c_doomhead[5467] = 5'h00;
assign _c_doomhead[5468] = 5'h00;
assign _c_doomhead[5469] = 5'h00;
assign _c_doomhead[5470] = 5'h00;
assign _c_doomhead[5471] = 5'h00;
assign _c_doomhead[5472] = 5'h00;
assign _c_doomhead[5473] = 5'h00;
assign _c_doomhead[5474] = 5'h00;
assign _c_doomhead[5475] = 5'h00;
assign _c_doomhead[5476] = 5'h11;
assign _c_doomhead[5477] = 5'h05;
assign _c_doomhead[5478] = 5'h06;
assign _c_doomhead[5479] = 5'h06;
assign _c_doomhead[5480] = 5'h1c;
assign _c_doomhead[5481] = 5'h1c;
assign _c_doomhead[5482] = 5'h0a;
assign _c_doomhead[5483] = 5'h0a;
assign _c_doomhead[5484] = 5'h03;
assign _c_doomhead[5485] = 5'h03;
assign _c_doomhead[5486] = 5'h08;
assign _c_doomhead[5487] = 5'h01;
assign _c_doomhead[5488] = 5'h03;
assign _c_doomhead[5489] = 5'h07;
assign _c_doomhead[5490] = 5'h09;
assign _c_doomhead[5491] = 5'h1b;
assign _c_doomhead[5492] = 5'h1b;
assign _c_doomhead[5493] = 5'h0a;
assign _c_doomhead[5494] = 5'h08;
assign _c_doomhead[5495] = 5'h07;
assign _c_doomhead[5496] = 5'h05;
assign _c_doomhead[5497] = 5'h11;
assign _c_doomhead[5498] = 5'h00;
assign _c_doomhead[5499] = 5'h00;
assign _c_doomhead[5500] = 5'h00;
assign _c_doomhead[5501] = 5'h00;
assign _c_doomhead[5502] = 5'h00;
assign _c_doomhead[5503] = 5'h00;
assign _c_doomhead[5504] = 5'h00;
assign _c_doomhead[5505] = 5'h00;
assign _c_doomhead[5506] = 5'h00;
assign _c_doomhead[5507] = 5'h0a;
assign _c_doomhead[5508] = 5'h17;
assign _c_doomhead[5509] = 5'h05;
assign _c_doomhead[5510] = 5'h01;
assign _c_doomhead[5511] = 5'h04;
assign _c_doomhead[5512] = 5'h1c;
assign _c_doomhead[5513] = 5'h1b;
assign _c_doomhead[5514] = 5'h0c;
assign _c_doomhead[5515] = 5'h18;
assign _c_doomhead[5516] = 5'h12;
assign _c_doomhead[5517] = 5'h03;
assign _c_doomhead[5518] = 5'h0a;
assign _c_doomhead[5519] = 5'h0a;
assign _c_doomhead[5520] = 5'h0c;
assign _c_doomhead[5521] = 5'h12;
assign _c_doomhead[5522] = 5'h14;
assign _c_doomhead[5523] = 5'h1b;
assign _c_doomhead[5524] = 5'h0e;
assign _c_doomhead[5525] = 5'h04;
assign _c_doomhead[5526] = 5'h04;
assign _c_doomhead[5527] = 5'h01;
assign _c_doomhead[5528] = 5'h05;
assign _c_doomhead[5529] = 5'h17;
assign _c_doomhead[5530] = 5'h0a;
assign _c_doomhead[5531] = 5'h00;
assign _c_doomhead[5532] = 5'h00;
assign _c_doomhead[5533] = 5'h00;
assign _c_doomhead[5534] = 5'h00;
assign _c_doomhead[5535] = 5'h00;
assign _c_doomhead[5536] = 5'h00;
assign _c_doomhead[5537] = 5'h00;
assign _c_doomhead[5538] = 5'h00;
assign _c_doomhead[5539] = 5'h0a;
assign _c_doomhead[5540] = 5'h04;
assign _c_doomhead[5541] = 5'h05;
assign _c_doomhead[5542] = 5'h06;
assign _c_doomhead[5543] = 5'h14;
assign _c_doomhead[5544] = 5'h1b;
assign _c_doomhead[5545] = 5'h1b;
assign _c_doomhead[5546] = 5'h10;
assign _c_doomhead[5547] = 5'h04;
assign _c_doomhead[5548] = 5'h08;
assign _c_doomhead[5549] = 5'h14;
assign _c_doomhead[5550] = 5'h12;
assign _c_doomhead[5551] = 5'h0c;
assign _c_doomhead[5552] = 5'h12;
assign _c_doomhead[5553] = 5'h0a;
assign _c_doomhead[5554] = 5'h04;
assign _c_doomhead[5555] = 5'h10;
assign _c_doomhead[5556] = 5'h01;
assign _c_doomhead[5557] = 5'h0b;
assign _c_doomhead[5558] = 5'h14;
assign _c_doomhead[5559] = 5'h06;
assign _c_doomhead[5560] = 5'h05;
assign _c_doomhead[5561] = 5'h04;
assign _c_doomhead[5562] = 5'h0a;
assign _c_doomhead[5563] = 5'h00;
assign _c_doomhead[5564] = 5'h00;
assign _c_doomhead[5565] = 5'h00;
assign _c_doomhead[5566] = 5'h00;
assign _c_doomhead[5567] = 5'h00;
assign _c_doomhead[5568] = 5'h00;
assign _c_doomhead[5569] = 5'h00;
assign _c_doomhead[5570] = 5'h00;
assign _c_doomhead[5571] = 5'h01;
assign _c_doomhead[5572] = 5'h04;
assign _c_doomhead[5573] = 5'h02;
assign _c_doomhead[5574] = 5'h04;
assign _c_doomhead[5575] = 5'h01;
assign _c_doomhead[5576] = 5'h17;
assign _c_doomhead[5577] = 5'h1d;
assign _c_doomhead[5578] = 5'h14;
assign _c_doomhead[5579] = 5'h10;
assign _c_doomhead[5580] = 5'h05;
assign _c_doomhead[5581] = 5'h01;
assign _c_doomhead[5582] = 5'h14;
assign _c_doomhead[5583] = 5'h0f;
assign _c_doomhead[5584] = 5'h01;
assign _c_doomhead[5585] = 5'h05;
assign _c_doomhead[5586] = 5'h10;
assign _c_doomhead[5587] = 5'h1d;
assign _c_doomhead[5588] = 5'h14;
assign _c_doomhead[5589] = 5'h17;
assign _c_doomhead[5590] = 5'h01;
assign _c_doomhead[5591] = 5'h04;
assign _c_doomhead[5592] = 5'h08;
assign _c_doomhead[5593] = 5'h04;
assign _c_doomhead[5594] = 5'h01;
assign _c_doomhead[5595] = 5'h00;
assign _c_doomhead[5596] = 5'h00;
assign _c_doomhead[5597] = 5'h00;
assign _c_doomhead[5598] = 5'h00;
assign _c_doomhead[5599] = 5'h00;
assign _c_doomhead[5600] = 5'h00;
assign _c_doomhead[5601] = 5'h00;
assign _c_doomhead[5602] = 5'h00;
assign _c_doomhead[5603] = 5'h04;
assign _c_doomhead[5604] = 5'h02;
assign _c_doomhead[5605] = 5'h02;
assign _c_doomhead[5606] = 5'h08;
assign _c_doomhead[5607] = 5'h0e;
assign _c_doomhead[5608] = 5'h1d;
assign _c_doomhead[5609] = 5'h05;
assign _c_doomhead[5610] = 5'h17;
assign _c_doomhead[5611] = 5'h14;
assign _c_doomhead[5612] = 5'h17;
assign _c_doomhead[5613] = 5'h0e;
assign _c_doomhead[5614] = 5'h09;
assign _c_doomhead[5615] = 5'h18;
assign _c_doomhead[5616] = 5'h0e;
assign _c_doomhead[5617] = 5'h17;
assign _c_doomhead[5618] = 5'h1d;
assign _c_doomhead[5619] = 5'h17;
assign _c_doomhead[5620] = 5'h05;
assign _c_doomhead[5621] = 5'h14;
assign _c_doomhead[5622] = 5'h0e;
assign _c_doomhead[5623] = 5'h08;
assign _c_doomhead[5624] = 5'h08;
assign _c_doomhead[5625] = 5'h02;
assign _c_doomhead[5626] = 5'h04;
assign _c_doomhead[5627] = 5'h00;
assign _c_doomhead[5628] = 5'h00;
assign _c_doomhead[5629] = 5'h00;
assign _c_doomhead[5630] = 5'h00;
assign _c_doomhead[5631] = 5'h00;
assign _c_doomhead[5632] = 5'h00;
assign _c_doomhead[5633] = 5'h00;
assign _c_doomhead[5634] = 5'h00;
assign _c_doomhead[5635] = 5'h08;
assign _c_doomhead[5636] = 5'h02;
assign _c_doomhead[5637] = 5'h08;
assign _c_doomhead[5638] = 5'h0c;
assign _c_doomhead[5639] = 5'h0a;
assign _c_doomhead[5640] = 5'h02;
assign _c_doomhead[5641] = 5'h1b;
assign _c_doomhead[5642] = 5'h1b;
assign _c_doomhead[5643] = 5'h0c;
assign _c_doomhead[5644] = 5'h18;
assign _c_doomhead[5645] = 5'h01;
assign _c_doomhead[5646] = 5'h0f;
assign _c_doomhead[5647] = 5'h12;
assign _c_doomhead[5648] = 5'h01;
assign _c_doomhead[5649] = 5'h18;
assign _c_doomhead[5650] = 5'h0c;
assign _c_doomhead[5651] = 5'h1b;
assign _c_doomhead[5652] = 5'h1b;
assign _c_doomhead[5653] = 5'h02;
assign _c_doomhead[5654] = 5'h0a;
assign _c_doomhead[5655] = 5'h0c;
assign _c_doomhead[5656] = 5'h08;
assign _c_doomhead[5657] = 5'h02;
assign _c_doomhead[5658] = 5'h08;
assign _c_doomhead[5659] = 5'h00;
assign _c_doomhead[5660] = 5'h00;
assign _c_doomhead[5661] = 5'h00;
assign _c_doomhead[5662] = 5'h00;
assign _c_doomhead[5663] = 5'h00;
assign _c_doomhead[5664] = 5'h00;
assign _c_doomhead[5665] = 5'h00;
assign _c_doomhead[5666] = 5'h00;
assign _c_doomhead[5667] = 5'h01;
assign _c_doomhead[5668] = 5'h02;
assign _c_doomhead[5669] = 5'h01;
assign _c_doomhead[5670] = 5'h0c;
assign _c_doomhead[5671] = 5'h12;
assign _c_doomhead[5672] = 5'h0d;
assign _c_doomhead[5673] = 5'h02;
assign _c_doomhead[5674] = 5'h08;
assign _c_doomhead[5675] = 5'h0c;
assign _c_doomhead[5676] = 5'h16;
assign _c_doomhead[5677] = 5'h0d;
assign _c_doomhead[5678] = 5'h0c;
assign _c_doomhead[5679] = 5'h18;
assign _c_doomhead[5680] = 5'h0d;
assign _c_doomhead[5681] = 5'h16;
assign _c_doomhead[5682] = 5'h0c;
assign _c_doomhead[5683] = 5'h08;
assign _c_doomhead[5684] = 5'h02;
assign _c_doomhead[5685] = 5'h0a;
assign _c_doomhead[5686] = 5'h12;
assign _c_doomhead[5687] = 5'h0c;
assign _c_doomhead[5688] = 5'h01;
assign _c_doomhead[5689] = 5'h02;
assign _c_doomhead[5690] = 5'h01;
assign _c_doomhead[5691] = 5'h00;
assign _c_doomhead[5692] = 5'h00;
assign _c_doomhead[5693] = 5'h00;
assign _c_doomhead[5694] = 5'h00;
assign _c_doomhead[5695] = 5'h00;
assign _c_doomhead[5696] = 5'h00;
assign _c_doomhead[5697] = 5'h00;
assign _c_doomhead[5698] = 5'h00;
assign _c_doomhead[5699] = 5'h00;
assign _c_doomhead[5700] = 5'h02;
assign _c_doomhead[5701] = 5'h01;
assign _c_doomhead[5702] = 5'h0f;
assign _c_doomhead[5703] = 5'h12;
assign _c_doomhead[5704] = 5'h0f;
assign _c_doomhead[5705] = 5'h0d;
assign _c_doomhead[5706] = 5'h16;
assign _c_doomhead[5707] = 5'h19;
assign _c_doomhead[5708] = 5'h18;
assign _c_doomhead[5709] = 5'h0d;
assign _c_doomhead[5710] = 5'h18;
assign _c_doomhead[5711] = 5'h16;
assign _c_doomhead[5712] = 5'h0d;
assign _c_doomhead[5713] = 5'h18;
assign _c_doomhead[5714] = 5'h18;
assign _c_doomhead[5715] = 5'h1e;
assign _c_doomhead[5716] = 5'h1e;
assign _c_doomhead[5717] = 5'h18;
assign _c_doomhead[5718] = 5'h12;
assign _c_doomhead[5719] = 5'h0f;
assign _c_doomhead[5720] = 5'h01;
assign _c_doomhead[5721] = 5'h02;
assign _c_doomhead[5722] = 5'h00;
assign _c_doomhead[5723] = 5'h00;
assign _c_doomhead[5724] = 5'h00;
assign _c_doomhead[5725] = 5'h00;
assign _c_doomhead[5726] = 5'h00;
assign _c_doomhead[5727] = 5'h00;
assign _c_doomhead[5728] = 5'h00;
assign _c_doomhead[5729] = 5'h00;
assign _c_doomhead[5730] = 5'h00;
assign _c_doomhead[5731] = 5'h00;
assign _c_doomhead[5732] = 5'h02;
assign _c_doomhead[5733] = 5'h01;
assign _c_doomhead[5734] = 5'h01;
assign _c_doomhead[5735] = 5'h0a;
assign _c_doomhead[5736] = 5'h1d;
assign _c_doomhead[5737] = 5'h12;
assign _c_doomhead[5738] = 5'h0c;
assign _c_doomhead[5739] = 5'h01;
assign _c_doomhead[5740] = 5'h0b;
assign _c_doomhead[5741] = 5'h07;
assign _c_doomhead[5742] = 5'h00;
assign _c_doomhead[5743] = 5'h00;
assign _c_doomhead[5744] = 5'h07;
assign _c_doomhead[5745] = 5'h0b;
assign _c_doomhead[5746] = 5'h01;
assign _c_doomhead[5747] = 5'h1e;
assign _c_doomhead[5748] = 5'h1e;
assign _c_doomhead[5749] = 5'h0b;
assign _c_doomhead[5750] = 5'h0f;
assign _c_doomhead[5751] = 5'h01;
assign _c_doomhead[5752] = 5'h01;
assign _c_doomhead[5753] = 5'h02;
assign _c_doomhead[5754] = 5'h00;
assign _c_doomhead[5755] = 5'h00;
assign _c_doomhead[5756] = 5'h00;
assign _c_doomhead[5757] = 5'h00;
assign _c_doomhead[5758] = 5'h00;
assign _c_doomhead[5759] = 5'h00;
assign _c_doomhead[5760] = 5'h00;
assign _c_doomhead[5761] = 5'h00;
assign _c_doomhead[5762] = 5'h00;
assign _c_doomhead[5763] = 5'h00;
assign _c_doomhead[5764] = 5'h02;
assign _c_doomhead[5765] = 5'h09;
assign _c_doomhead[5766] = 5'h15;
assign _c_doomhead[5767] = 5'h1d;
assign _c_doomhead[5768] = 5'h09;
assign _c_doomhead[5769] = 5'h12;
assign _c_doomhead[5770] = 5'h01;
assign _c_doomhead[5771] = 5'h08;
assign _c_doomhead[5772] = 5'h0e;
assign _c_doomhead[5773] = 5'h06;
assign _c_doomhead[5774] = 5'h08;
assign _c_doomhead[5775] = 5'h08;
assign _c_doomhead[5776] = 5'h06;
assign _c_doomhead[5777] = 5'h0e;
assign _c_doomhead[5778] = 5'h08;
assign _c_doomhead[5779] = 5'h1e;
assign _c_doomhead[5780] = 5'h1a;
assign _c_doomhead[5781] = 5'h09;
assign _c_doomhead[5782] = 5'h15;
assign _c_doomhead[5783] = 5'h15;
assign _c_doomhead[5784] = 5'h09;
assign _c_doomhead[5785] = 5'h02;
assign _c_doomhead[5786] = 5'h00;
assign _c_doomhead[5787] = 5'h00;
assign _c_doomhead[5788] = 5'h00;
assign _c_doomhead[5789] = 5'h00;
assign _c_doomhead[5790] = 5'h00;
assign _c_doomhead[5791] = 5'h00;
assign _c_doomhead[5792] = 5'h00;
assign _c_doomhead[5793] = 5'h00;
assign _c_doomhead[5794] = 5'h00;
assign _c_doomhead[5795] = 5'h00;
assign _c_doomhead[5796] = 5'h00;
assign _c_doomhead[5797] = 5'h01;
assign _c_doomhead[5798] = 5'h01;
assign _c_doomhead[5799] = 5'h1d;
assign _c_doomhead[5800] = 5'h09;
assign _c_doomhead[5801] = 5'h0d;
assign _c_doomhead[5802] = 5'h04;
assign _c_doomhead[5803] = 5'h0a;
assign _c_doomhead[5804] = 5'h1d;
assign _c_doomhead[5805] = 5'h1a;
assign _c_doomhead[5806] = 5'h04;
assign _c_doomhead[5807] = 5'h04;
assign _c_doomhead[5808] = 5'h1a;
assign _c_doomhead[5809] = 5'h1d;
assign _c_doomhead[5810] = 5'h0a;
assign _c_doomhead[5811] = 5'h04;
assign _c_doomhead[5812] = 5'h1a;
assign _c_doomhead[5813] = 5'h09;
assign _c_doomhead[5814] = 5'h08;
assign _c_doomhead[5815] = 5'h09;
assign _c_doomhead[5816] = 5'h01;
assign _c_doomhead[5817] = 5'h00;
assign _c_doomhead[5818] = 5'h00;
assign _c_doomhead[5819] = 5'h00;
assign _c_doomhead[5820] = 5'h00;
assign _c_doomhead[5821] = 5'h00;
assign _c_doomhead[5822] = 5'h00;
assign _c_doomhead[5823] = 5'h00;
assign _c_doomhead[5824] = 5'h00;
assign _c_doomhead[5825] = 5'h00;
assign _c_doomhead[5826] = 5'h00;
assign _c_doomhead[5827] = 5'h00;
assign _c_doomhead[5828] = 5'h00;
assign _c_doomhead[5829] = 5'h15;
assign _c_doomhead[5830] = 5'h09;
assign _c_doomhead[5831] = 5'h15;
assign _c_doomhead[5832] = 5'h1b;
assign _c_doomhead[5833] = 5'h0c;
assign _c_doomhead[5834] = 5'h06;
assign _c_doomhead[5835] = 5'h0a;
assign _c_doomhead[5836] = 5'h1c;
assign _c_doomhead[5837] = 5'h1a;
assign _c_doomhead[5838] = 5'h1c;
assign _c_doomhead[5839] = 5'h1c;
assign _c_doomhead[5840] = 5'h1a;
assign _c_doomhead[5841] = 5'h1b;
assign _c_doomhead[5842] = 5'h0a;
assign _c_doomhead[5843] = 5'h06;
assign _c_doomhead[5844] = 5'h1a;
assign _c_doomhead[5845] = 5'h09;
assign _c_doomhead[5846] = 5'h15;
assign _c_doomhead[5847] = 5'h0f;
assign _c_doomhead[5848] = 5'h15;
assign _c_doomhead[5849] = 5'h00;
assign _c_doomhead[5850] = 5'h00;
assign _c_doomhead[5851] = 5'h00;
assign _c_doomhead[5852] = 5'h00;
assign _c_doomhead[5853] = 5'h00;
assign _c_doomhead[5854] = 5'h00;
assign _c_doomhead[5855] = 5'h00;
assign _c_doomhead[5856] = 5'h00;
assign _c_doomhead[5857] = 5'h00;
assign _c_doomhead[5858] = 5'h00;
assign _c_doomhead[5859] = 5'h00;
assign _c_doomhead[5860] = 5'h00;
assign _c_doomhead[5861] = 5'h00;
assign _c_doomhead[5862] = 5'h01;
assign _c_doomhead[5863] = 5'h15;
assign _c_doomhead[5864] = 5'h1b;
assign _c_doomhead[5865] = 5'h0f;
assign _c_doomhead[5866] = 5'h07;
assign _c_doomhead[5867] = 5'h0d;
assign _c_doomhead[5868] = 5'h1a;
assign _c_doomhead[5869] = 5'h1a;
assign _c_doomhead[5870] = 5'h06;
assign _c_doomhead[5871] = 5'h06;
assign _c_doomhead[5872] = 5'h1a;
assign _c_doomhead[5873] = 5'h1c;
assign _c_doomhead[5874] = 5'h0f;
assign _c_doomhead[5875] = 5'h07;
assign _c_doomhead[5876] = 5'h1c;
assign _c_doomhead[5877] = 5'h07;
assign _c_doomhead[5878] = 5'h15;
assign _c_doomhead[5879] = 5'h09;
assign _c_doomhead[5880] = 5'h00;
assign _c_doomhead[5881] = 5'h00;
assign _c_doomhead[5882] = 5'h00;
assign _c_doomhead[5883] = 5'h00;
assign _c_doomhead[5884] = 5'h00;
assign _c_doomhead[5885] = 5'h00;
assign _c_doomhead[5886] = 5'h00;
assign _c_doomhead[5887] = 5'h00;
assign _c_doomhead[5888] = 5'h00;
assign _c_doomhead[5889] = 5'h00;
assign _c_doomhead[5890] = 5'h00;
assign _c_doomhead[5891] = 5'h00;
assign _c_doomhead[5892] = 5'h00;
assign _c_doomhead[5893] = 5'h00;
assign _c_doomhead[5894] = 5'h08;
assign _c_doomhead[5895] = 5'h15;
assign _c_doomhead[5896] = 5'h1b;
assign _c_doomhead[5897] = 5'h0f;
assign _c_doomhead[5898] = 5'h07;
assign _c_doomhead[5899] = 5'h0a;
assign _c_doomhead[5900] = 5'h1c;
assign _c_doomhead[5901] = 5'h1c;
assign _c_doomhead[5902] = 5'h1a;
assign _c_doomhead[5903] = 5'h1a;
assign _c_doomhead[5904] = 5'h1c;
assign _c_doomhead[5905] = 5'h1c;
assign _c_doomhead[5906] = 5'h1e;
assign _c_doomhead[5907] = 5'h07;
assign _c_doomhead[5908] = 5'h1c;
assign _c_doomhead[5909] = 5'h08;
assign _c_doomhead[5910] = 5'h15;
assign _c_doomhead[5911] = 5'h08;
assign _c_doomhead[5912] = 5'h00;
assign _c_doomhead[5913] = 5'h00;
assign _c_doomhead[5914] = 5'h00;
assign _c_doomhead[5915] = 5'h00;
assign _c_doomhead[5916] = 5'h00;
assign _c_doomhead[5917] = 5'h00;
assign _c_doomhead[5918] = 5'h00;
assign _c_doomhead[5919] = 5'h00;
assign _c_doomhead[5920] = 5'h00;
assign _c_doomhead[5921] = 5'h00;
assign _c_doomhead[5922] = 5'h00;
assign _c_doomhead[5923] = 5'h00;
assign _c_doomhead[5924] = 5'h00;
assign _c_doomhead[5925] = 5'h00;
assign _c_doomhead[5926] = 5'h06;
assign _c_doomhead[5927] = 5'h15;
assign _c_doomhead[5928] = 5'h1a;
assign _c_doomhead[5929] = 5'h09;
assign _c_doomhead[5930] = 5'h0b;
assign _c_doomhead[5931] = 5'h07;
assign _c_doomhead[5932] = 5'h1c;
assign _c_doomhead[5933] = 5'h17;
assign _c_doomhead[5934] = 5'h17;
assign _c_doomhead[5935] = 5'h17;
assign _c_doomhead[5936] = 5'h17;
assign _c_doomhead[5937] = 5'h1c;
assign _c_doomhead[5938] = 5'h1e;
assign _c_doomhead[5939] = 5'h1a;
assign _c_doomhead[5940] = 5'h1c;
assign _c_doomhead[5941] = 5'h06;
assign _c_doomhead[5942] = 5'h15;
assign _c_doomhead[5943] = 5'h06;
assign _c_doomhead[5944] = 5'h00;
assign _c_doomhead[5945] = 5'h00;
assign _c_doomhead[5946] = 5'h00;
assign _c_doomhead[5947] = 5'h00;
assign _c_doomhead[5948] = 5'h00;
assign _c_doomhead[5949] = 5'h00;
assign _c_doomhead[5950] = 5'h00;
assign _c_doomhead[5951] = 5'h00;
assign _c_doomhead[5952] = 5'h00;
assign _c_doomhead[5953] = 5'h00;
assign _c_doomhead[5954] = 5'h00;
assign _c_doomhead[5955] = 5'h00;
assign _c_doomhead[5956] = 5'h00;
assign _c_doomhead[5957] = 5'h00;
assign _c_doomhead[5958] = 5'h00;
assign _c_doomhead[5959] = 5'h15;
assign _c_doomhead[5960] = 5'h1c;
assign _c_doomhead[5961] = 5'h01;
assign _c_doomhead[5962] = 5'h0f;
assign _c_doomhead[5963] = 5'h08;
assign _c_doomhead[5964] = 5'h1b;
assign _c_doomhead[5965] = 5'h1c;
assign _c_doomhead[5966] = 5'h17;
assign _c_doomhead[5967] = 5'h17;
assign _c_doomhead[5968] = 5'h1c;
assign _c_doomhead[5969] = 5'h1c;
assign _c_doomhead[5970] = 5'h1e;
assign _c_doomhead[5971] = 5'h1a;
assign _c_doomhead[5972] = 5'h1a;
assign _c_doomhead[5973] = 5'h06;
assign _c_doomhead[5974] = 5'h15;
assign _c_doomhead[5975] = 5'h00;
assign _c_doomhead[5976] = 5'h00;
assign _c_doomhead[5977] = 5'h00;
assign _c_doomhead[5978] = 5'h00;
assign _c_doomhead[5979] = 5'h00;
assign _c_doomhead[5980] = 5'h00;
assign _c_doomhead[5981] = 5'h00;
assign _c_doomhead[5982] = 5'h00;
assign _c_doomhead[5983] = 5'h00;
assign _c_doomhead[5984] = 5'h00;
assign _c_doomhead[5985] = 5'h00;
assign _c_doomhead[5986] = 5'h00;
assign _c_doomhead[5987] = 5'h00;
assign _c_doomhead[5988] = 5'h00;
assign _c_doomhead[5989] = 5'h00;
assign _c_doomhead[5990] = 5'h00;
assign _c_doomhead[5991] = 5'h06;
assign _c_doomhead[5992] = 5'h1c;
assign _c_doomhead[5993] = 5'h08;
assign _c_doomhead[5994] = 5'h0c;
assign _c_doomhead[5995] = 5'h09;
assign _c_doomhead[5996] = 5'h1a;
assign _c_doomhead[5997] = 5'h1d;
assign _c_doomhead[5998] = 5'h1e;
assign _c_doomhead[5999] = 5'h1e;
assign _c_doomhead[6000] = 5'h1d;
assign _c_doomhead[6001] = 5'h1a;
assign _c_doomhead[6002] = 5'h0f;
assign _c_doomhead[6003] = 5'h0c;
assign _c_doomhead[6004] = 5'h1a;
assign _c_doomhead[6005] = 5'h06;
assign _c_doomhead[6006] = 5'h06;
assign _c_doomhead[6007] = 5'h00;
assign _c_doomhead[6008] = 5'h00;
assign _c_doomhead[6009] = 5'h00;
assign _c_doomhead[6010] = 5'h00;
assign _c_doomhead[6011] = 5'h00;
assign _c_doomhead[6012] = 5'h00;
assign _c_doomhead[6013] = 5'h00;
assign _c_doomhead[6014] = 5'h00;
assign _c_doomhead[6015] = 5'h00;
assign _c_doomhead[6016] = 5'h00;
assign _c_doomhead[6017] = 5'h00;
assign _c_doomhead[6018] = 5'h00;
assign _c_doomhead[6019] = 5'h00;
assign _c_doomhead[6020] = 5'h00;
assign _c_doomhead[6021] = 5'h00;
assign _c_doomhead[6022] = 5'h00;
assign _c_doomhead[6023] = 5'h00;
assign _c_doomhead[6024] = 5'h1c;
assign _c_doomhead[6025] = 5'h15;
assign _c_doomhead[6026] = 5'h0a;
assign _c_doomhead[6027] = 5'h0b;
assign _c_doomhead[6028] = 5'h1c;
assign _c_doomhead[6029] = 5'h1c;
assign _c_doomhead[6030] = 5'h1d;
assign _c_doomhead[6031] = 5'h1d;
assign _c_doomhead[6032] = 5'h1a;
assign _c_doomhead[6033] = 5'h1c;
assign _c_doomhead[6034] = 5'h0b;
assign _c_doomhead[6035] = 5'h0a;
assign _c_doomhead[6036] = 5'h1c;
assign _c_doomhead[6037] = 5'h06;
assign _c_doomhead[6038] = 5'h00;
assign _c_doomhead[6039] = 5'h00;
assign _c_doomhead[6040] = 5'h00;
assign _c_doomhead[6041] = 5'h00;
assign _c_doomhead[6042] = 5'h00;
assign _c_doomhead[6043] = 5'h00;
assign _c_doomhead[6044] = 5'h00;
assign _c_doomhead[6045] = 5'h00;
assign _c_doomhead[6046] = 5'h00;
assign _c_doomhead[6047] = 5'h00;
assign _c_doomhead[6048] = 5'h00;
assign _c_doomhead[6049] = 5'h00;
assign _c_doomhead[6050] = 5'h00;
assign _c_doomhead[6051] = 5'h00;
assign _c_doomhead[6052] = 5'h00;
assign _c_doomhead[6053] = 5'h00;
assign _c_doomhead[6054] = 5'h00;
assign _c_doomhead[6055] = 5'h00;
assign _c_doomhead[6056] = 5'h00;
assign _c_doomhead[6057] = 5'h1c;
assign _c_doomhead[6058] = 5'h01;
assign _c_doomhead[6059] = 5'h0b;
assign _c_doomhead[6060] = 5'h1c;
assign _c_doomhead[6061] = 5'h1c;
assign _c_doomhead[6062] = 5'h15;
assign _c_doomhead[6063] = 5'h15;
assign _c_doomhead[6064] = 5'h1a;
assign _c_doomhead[6065] = 5'h1c;
assign _c_doomhead[6066] = 5'h0b;
assign _c_doomhead[6067] = 5'h01;
assign _c_doomhead[6068] = 5'h1c;
assign _c_doomhead[6069] = 5'h00;
assign _c_doomhead[6070] = 5'h00;
assign _c_doomhead[6071] = 5'h00;
assign _c_doomhead[6072] = 5'h00;
assign _c_doomhead[6073] = 5'h00;
assign _c_doomhead[6074] = 5'h00;
assign _c_doomhead[6075] = 5'h00;
assign _c_doomhead[6076] = 5'h00;
assign _c_doomhead[6077] = 5'h00;
assign _c_doomhead[6078] = 5'h00;
assign _c_doomhead[6079] = 5'h00;
assign _c_doomhead[6080] = 5'h00;
assign _c_doomhead[6081] = 5'h00;
assign _c_doomhead[6082] = 5'h00;
assign _c_doomhead[6083] = 5'h00;
assign _c_doomhead[6084] = 5'h00;
assign _c_doomhead[6085] = 5'h00;
assign _c_doomhead[6086] = 5'h00;
assign _c_doomhead[6087] = 5'h00;
assign _c_doomhead[6088] = 5'h00;
assign _c_doomhead[6089] = 5'h00;
assign _c_doomhead[6090] = 5'h06;
assign _c_doomhead[6091] = 5'h07;
assign _c_doomhead[6092] = 5'h03;
assign _c_doomhead[6093] = 5'h1c;
assign _c_doomhead[6094] = 5'h1e;
assign _c_doomhead[6095] = 5'h1e;
assign _c_doomhead[6096] = 5'h1e;
assign _c_doomhead[6097] = 5'h1c;
assign _c_doomhead[6098] = 5'h07;
assign _c_doomhead[6099] = 5'h1a;
assign _c_doomhead[6100] = 5'h00;
assign _c_doomhead[6101] = 5'h00;
assign _c_doomhead[6102] = 5'h00;
assign _c_doomhead[6103] = 5'h00;
assign _c_doomhead[6104] = 5'h00;
assign _c_doomhead[6105] = 5'h00;
assign _c_doomhead[6106] = 5'h00;
assign _c_doomhead[6107] = 5'h00;
assign _c_doomhead[6108] = 5'h00;
assign _c_doomhead[6109] = 5'h00;
assign _c_doomhead[6110] = 5'h00;
assign _c_doomhead[6111] = 5'h00;
assign _c_doomhead[6112] = 5'h00;
assign _c_doomhead[6113] = 5'h00;
assign _c_doomhead[6114] = 5'h00;
assign _c_doomhead[6115] = 5'h00;
assign _c_doomhead[6116] = 5'h00;
assign _c_doomhead[6117] = 5'h00;
assign _c_doomhead[6118] = 5'h00;
assign _c_doomhead[6119] = 5'h00;
assign _c_doomhead[6120] = 5'h00;
assign _c_doomhead[6121] = 5'h00;
assign _c_doomhead[6122] = 5'h00;
assign _c_doomhead[6123] = 5'h00;
assign _c_doomhead[6124] = 5'h00;
assign _c_doomhead[6125] = 5'h00;
assign _c_doomhead[6126] = 5'h00;
assign _c_doomhead[6127] = 5'h00;
assign _c_doomhead[6128] = 5'h00;
assign _c_doomhead[6129] = 5'h00;
assign _c_doomhead[6130] = 5'h00;
assign _c_doomhead[6131] = 5'h00;
assign _c_doomhead[6132] = 5'h00;
assign _c_doomhead[6133] = 5'h00;
assign _c_doomhead[6134] = 5'h00;
assign _c_doomhead[6135] = 5'h00;
assign _c_doomhead[6136] = 5'h00;
assign _c_doomhead[6137] = 5'h00;
assign _c_doomhead[6138] = 5'h00;
assign _c_doomhead[6139] = 5'h00;
assign _c_doomhead[6140] = 5'h00;
assign _c_doomhead[6141] = 5'h00;
assign _c_doomhead[6142] = 5'h00;
assign _c_doomhead[6143] = 5'h00;
wire  [23:0] _c_sub666[31:0];
assign _c_sub666[0] = 169626;
assign _c_sub666[1] = 144845;
assign _c_sub666[2] = 95240;
assign _c_sub666[3] = 49796;
assign _c_sub666[4] = 107593;
assign _c_sub666[5] = 74566;
assign _c_sub666[6] = 120010;
assign _c_sub666[7] = 157198;
assign _c_sub666[8] = 136524;
assign _c_sub666[9] = 165519;
assign _c_sub666[10] = 182033;
assign _c_sub666[11] = 173776;
assign _c_sub666[12] = 210964;
assign _c_sub666[13] = 219286;
assign _c_sub666[14] = 82887;
assign _c_sub666[15] = 194450;
assign _c_sub666[16] = 62149;
assign _c_sub666[17] = 41475;
assign _c_sub666[18] = 235930;
assign _c_sub666[19] = 206803;
assign _c_sub666[20] = 227608;
assign _c_sub666[21] = 128267;
assign _c_sub666[22] = 261028;
assign _c_sub666[23] = 0;
assign _c_sub666[24] = 252574;
assign _c_sub666[25] = 244252;
assign _c_sub666[26] = 144010;
assign _c_sub666[27] = 152267;
assign _c_sub666[28] = 127366;
assign _c_sub666[29] = 168911;
assign _c_sub666[30] = 177233;
assign _c_sub666[31] = 157060;
// ===============

always @(posedge clock) begin
end

endmodule


module M_main (
in_ui,
out_uo,
inout_uio_oe,
inout_uio_i,
inout_uio_o,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [7:0] in_ui;
output  [7:0] out_uo;
output  [7:0] inout_uio_oe;
input  [7:0] inout_uio_i;
output  [7:0] inout_uio_o;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [1:0] _w_demo_video_r;
wire  [1:0] _w_demo_video_g;
wire  [1:0] _w_demo_video_b;
wire  [0:0] _w_demo_video_hs;
wire  [0:0] _w_demo_video_vs;

reg  [7:0] _d_uio_oenable;
reg  [7:0] _q_uio_oenable;
reg  [7:0] _d_uo;
reg  [7:0] _q_uo;
assign out_uo = _q_uo;
assign out_done = 0;
M_vga_demo_M_main_demo demo (
.out_video_r(_w_demo_video_r),
.out_video_g(_w_demo_video_g),
.out_video_b(_w_demo_video_b),
.out_video_hs(_w_demo_video_hs),
.out_video_vs(_w_demo_video_vs),
.reset(reset),
.clock(clock));


assign inout_uio_oe[0] = _q_uio_oenable[0];
assign inout_uio_o[0] = 1'b0;
assign inout_uio_oe[1] = _q_uio_oenable[1];
assign inout_uio_o[1] = 1'b0;
assign inout_uio_oe[2] = _q_uio_oenable[2];
assign inout_uio_o[2] = 1'b0;
assign inout_uio_oe[3] = _q_uio_oenable[3];
assign inout_uio_o[3] = 1'b0;
assign inout_uio_oe[4] = _q_uio_oenable[4];
assign inout_uio_o[4] = 1'b0;
assign inout_uio_oe[5] = _q_uio_oenable[5];
assign inout_uio_o[5] = 1'b0;
assign inout_uio_oe[6] = _q_uio_oenable[6];
assign inout_uio_o[6] = 1'b0;
assign inout_uio_oe[7] = _q_uio_oenable[7];
assign inout_uio_o[7] = 1'b0;

`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
_d_uio_oenable = _q_uio_oenable;
_d_uo = _q_uo;
// _always_pre
// __block_1
_d_uo[7+:1] = _w_demo_video_hs;

_d_uo[3+:1] = _w_demo_video_vs;

_d_uo[4+:1] = _w_demo_video_r[0+:1];

_d_uo[0+:1] = _w_demo_video_r[1+:1];

_d_uo[5+:1] = _w_demo_video_g[0+:1];

_d_uo[1+:1] = _w_demo_video_g[1+:1];

_d_uo[6+:1] = _w_demo_video_b[0+:1];

_d_uo[2+:1] = _w_demo_video_b[1+:1];

_d_uio_oenable = 8'b0;

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
_q_uio_oenable <= _d_uio_oenable;
_q_uo <= _d_uo;
end

endmodule
